--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_efdf1b1b05926829.vhd when simulating
-- the core, dmg_72_efdf1b1b05926829. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_efdf1b1b05926829 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_efdf1b1b05926829;

ARCHITECTURE dmg_72_efdf1b1b05926829_a OF dmg_72_efdf1b1b05926829 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_efdf1b1b05926829
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_efdf1b1b05926829 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_efdf1b1b05926829.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_efdf1b1b05926829
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_efdf1b1b05926829_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_ed810b6704650710.vhd when simulating
-- the core, cntr_11_0_ed810b6704650710. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_ed810b6704650710 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END cntr_11_0_ed810b6704650710;

ARCHITECTURE cntr_11_0_ed810b6704650710_a OF cntr_11_0_ed810b6704650710 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_ed810b6704650710
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_ed810b6704650710 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 12,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_ed810b6704650710
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_ed810b6704650710_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_53d3a85261e207bb.vhd when simulating
-- the core, bmg_72_53d3a85261e207bb. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_53d3a85261e207bb IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_53d3a85261e207bb;

ARCHITECTURE bmg_72_53d3a85261e207bb_a OF bmg_72_53d3a85261e207bb IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_53d3a85261e207bb
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_53d3a85261e207bb USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_53d3a85261e207bb.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_53d3a85261e207bb
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_53d3a85261e207bb_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_2f7113c203379501.vhd when simulating
-- the core, cntr_11_0_2f7113c203379501. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_2f7113c203379501 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
  );
END cntr_11_0_2f7113c203379501;

ARCHITECTURE cntr_11_0_2f7113c203379501_a OF cntr_11_0_2f7113c203379501 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_2f7113c203379501
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_2f7113c203379501 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 11,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_2f7113c203379501
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_2f7113c203379501_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_9f585cf1e3329833.vhd when simulating
-- the core, bmg_72_9f585cf1e3329833. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_9f585cf1e3329833 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_9f585cf1e3329833;

ARCHITECTURE bmg_72_9f585cf1e3329833_a OF bmg_72_9f585cf1e3329833 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_9f585cf1e3329833
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_9f585cf1e3329833 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 10,
      c_addrb_width => 10,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_9f585cf1e3329833.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 1024,
      c_read_depth_b => 1024,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 1024,
      c_write_depth_b => 1024,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_9f585cf1e3329833
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_9f585cf1e3329833_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_efa60dbe2ed9d35a.vhd when simulating
-- the core, cntr_11_0_efa60dbe2ed9d35a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_efa60dbe2ed9d35a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END cntr_11_0_efa60dbe2ed9d35a;

ARCHITECTURE cntr_11_0_efa60dbe2ed9d35a_a OF cntr_11_0_efa60dbe2ed9d35a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_efa60dbe2ed9d35a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_efa60dbe2ed9d35a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 3,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_efa60dbe2ed9d35a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_efa60dbe2ed9d35a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_796a9d3dfbc0c498.vhd when simulating
-- the core, cntr_11_0_796a9d3dfbc0c498. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_796a9d3dfbc0c498 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END cntr_11_0_796a9d3dfbc0c498;

ARCHITECTURE cntr_11_0_796a9d3dfbc0c498_a OF cntr_11_0_796a9d3dfbc0c498 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_796a9d3dfbc0c498
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_796a9d3dfbc0c498 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_796a9d3dfbc0c498
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_796a9d3dfbc0c498_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_125dc8e6a3ba8cad.vhd when simulating
-- the core, cntr_11_0_125dc8e6a3ba8cad. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_125dc8e6a3ba8cad IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END cntr_11_0_125dc8e6a3ba8cad;

ARCHITECTURE cntr_11_0_125dc8e6a3ba8cad_a OF cntr_11_0_125dc8e6a3ba8cad IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_125dc8e6a3ba8cad
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_125dc8e6a3ba8cad USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 13,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_125dc8e6a3ba8cad
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_125dc8e6a3ba8cad_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_a0497faccc62b6b2.vhd when simulating
-- the core, addsb_11_0_a0497faccc62b6b2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_a0497faccc62b6b2 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END addsb_11_0_a0497faccc62b6b2;

ARCHITECTURE addsb_11_0_a0497faccc62b6b2_a OF addsb_11_0_a0497faccc62b6b2 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_a0497faccc62b6b2
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_a0497faccc62b6b2 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 20,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000",
      c_b_width => 20,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 20,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_a0497faccc62b6b2
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_a0497faccc62b6b2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_d60ecc44fc05ecdd.vhd when simulating
-- the core, cntr_11_0_d60ecc44fc05ecdd. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_d60ecc44fc05ecdd IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END cntr_11_0_d60ecc44fc05ecdd;

ARCHITECTURE cntr_11_0_d60ecc44fc05ecdd_a OF cntr_11_0_d60ecc44fc05ecdd IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_d60ecc44fc05ecdd
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_d60ecc44fc05ecdd USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 6,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_d60ecc44fc05ecdd
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_d60ecc44fc05ecdd_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_ee60311bb9d0db53.vhd when simulating
-- the core, cntr_11_0_ee60311bb9d0db53. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_ee60311bb9d0db53 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END cntr_11_0_ee60311bb9d0db53;

ARCHITECTURE cntr_11_0_ee60311bb9d0db53_a OF cntr_11_0_ee60311bb9d0db53 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_ee60311bb9d0db53
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_ee60311bb9d0db53 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 5,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_ee60311bb9d0db53
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_ee60311bb9d0db53_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_756e5f183b33a31a.vhd when simulating
-- the core, bmg_72_756e5f183b33a31a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_756e5f183b33a31a IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_756e5f183b33a31a;

ARCHITECTURE bmg_72_756e5f183b33a31a_a OF bmg_72_756e5f183b33a31a IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_756e5f183b33a31a
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_756e5f183b33a31a USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 10,
      c_addrb_width => 10,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_756e5f183b33a31a.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 1024,
      c_read_depth_b => 1024,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 1024,
      c_write_depth_b => 1024,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_756e5f183b33a31a
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_756e5f183b33a31a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_3a3ea2f70b8548a5.vhd when simulating
-- the core, cntr_11_0_3a3ea2f70b8548a5. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_3a3ea2f70b8548a5 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END cntr_11_0_3a3ea2f70b8548a5;

ARCHITECTURE cntr_11_0_3a3ea2f70b8548a5_a OF cntr_11_0_3a3ea2f70b8548a5 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_3a3ea2f70b8548a5
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_3a3ea2f70b8548a5 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 3,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_3a3ea2f70b8548a5
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_3a3ea2f70b8548a5_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_461fd5d45cff2f9b.vhd when simulating
-- the core, cntr_11_0_461fd5d45cff2f9b. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_461fd5d45cff2f9b IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END cntr_11_0_461fd5d45cff2f9b;

ARCHITECTURE cntr_11_0_461fd5d45cff2f9b_a OF cntr_11_0_461fd5d45cff2f9b IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_461fd5d45cff2f9b
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_461fd5d45cff2f9b USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 13,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_461fd5d45cff2f9b
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_461fd5d45cff2f9b_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_99383d874600f8be.vhd when simulating
-- the core, cntr_11_0_99383d874600f8be. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_99383d874600f8be IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END cntr_11_0_99383d874600f8be;

ARCHITECTURE cntr_11_0_99383d874600f8be_a OF cntr_11_0_99383d874600f8be IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_99383d874600f8be
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_99383d874600f8be USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 2,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_99383d874600f8be
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_99383d874600f8be_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_87bb354a843dab37.vhd when simulating
-- the core, bmg_72_87bb354a843dab37. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_87bb354a843dab37 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_87bb354a843dab37;

ARCHITECTURE bmg_72_87bb354a843dab37_a OF bmg_72_87bb354a843dab37 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_87bb354a843dab37
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_87bb354a843dab37 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 8,
      c_addrb_width => 8,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_87bb354a843dab37.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 256,
      c_read_depth_b => 256,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 256,
      c_write_depth_b => 256,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_87bb354a843dab37
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_87bb354a843dab37_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_133a8817831fb97a.vhd when simulating
-- the core, cntr_11_0_133a8817831fb97a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_133a8817831fb97a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_133a8817831fb97a;

ARCHITECTURE cntr_11_0_133a8817831fb97a_a OF cntr_11_0_133a8817831fb97a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_133a8817831fb97a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_133a8817831fb97a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_133a8817831fb97a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_133a8817831fb97a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_b5cea772b1c370b5.vhd when simulating
-- the core, dmg_72_b5cea772b1c370b5. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_b5cea772b1c370b5 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END dmg_72_b5cea772b1c370b5;

ARCHITECTURE dmg_72_b5cea772b1c370b5_a OF dmg_72_b5cea772b1c370b5 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_b5cea772b1c370b5
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_b5cea772b1c370b5 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 12,
      c_default_data => "0",
      c_depth => 4096,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_b5cea772b1c370b5.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 12
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_b5cea772b1c370b5
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_b5cea772b1c370b5_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_59920783799a8e86.vhd when simulating
-- the core, addsb_11_0_59920783799a8e86. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_59920783799a8e86 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_59920783799a8e86;

ARCHITECTURE addsb_11_0_59920783799a8e86_a OF addsb_11_0_59920783799a8e86 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_59920783799a8e86
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_59920783799a8e86 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_59920783799a8e86
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_59920783799a8e86_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_cb1ffe90ceffe54f.vhd when simulating
-- the core, cntr_11_0_cb1ffe90ceffe54f. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_cb1ffe90ceffe54f IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END cntr_11_0_cb1ffe90ceffe54f;

ARCHITECTURE cntr_11_0_cb1ffe90ceffe54f_a OF cntr_11_0_cb1ffe90ceffe54f IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_cb1ffe90ceffe54f
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_cb1ffe90ceffe54f USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 6,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_cb1ffe90ceffe54f
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_cb1ffe90ceffe54f_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_08915946f5ebdf9c.vhd when simulating
-- the core, dmg_72_08915946f5ebdf9c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_08915946f5ebdf9c IS
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END dmg_72_08915946f5ebdf9c;

ARCHITECTURE dmg_72_08915946f5ebdf9c_a OF dmg_72_08915946f5ebdf9c IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_08915946f5ebdf9c
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_08915946f5ebdf9c USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 12,
      c_default_data => "0",
      c_depth => 4096,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_08915946f5ebdf9c.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 12
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_08915946f5ebdf9c
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_08915946f5ebdf9c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_a2916e7e77833dd6.vhd when simulating
-- the core, cntr_11_0_a2916e7e77833dd6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_a2916e7e77833dd6 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END cntr_11_0_a2916e7e77833dd6;

ARCHITECTURE cntr_11_0_a2916e7e77833dd6_a OF cntr_11_0_a2916e7e77833dd6 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_a2916e7e77833dd6
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_a2916e7e77833dd6 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 12,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_a2916e7e77833dd6
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_a2916e7e77833dd6_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_59143b4ed22b761d.vhd when simulating
-- the core, bmg_72_59143b4ed22b761d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_59143b4ed22b761d IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_59143b4ed22b761d;

ARCHITECTURE bmg_72_59143b4ed22b761d_a OF bmg_72_59143b4ed22b761d IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_59143b4ed22b761d
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_59143b4ed22b761d USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_59143b4ed22b761d.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 64,
      c_read_depth_b => 64,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 64,
      c_write_depth_b => 64,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_59143b4ed22b761d
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_59143b4ed22b761d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_c1a8b20e2e422729.vhd when simulating
-- the core, bmg_72_c1a8b20e2e422729. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_c1a8b20e2e422729 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_c1a8b20e2e422729;

ARCHITECTURE bmg_72_c1a8b20e2e422729_a OF bmg_72_c1a8b20e2e422729 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_c1a8b20e2e422729
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_c1a8b20e2e422729 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 9,
      c_addrb_width => 9,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_c1a8b20e2e422729.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 512,
      c_read_depth_b => 512,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 512,
      c_write_depth_b => 512,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_c1a8b20e2e422729
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_c1a8b20e2e422729_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_d5eedfa744d4da30.vhd when simulating
-- the core, cntr_11_0_d5eedfa744d4da30. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_d5eedfa744d4da30 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END cntr_11_0_d5eedfa744d4da30;

ARCHITECTURE cntr_11_0_d5eedfa744d4da30_a OF cntr_11_0_d5eedfa744d4da30 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_d5eedfa744d4da30
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_d5eedfa744d4da30 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 5,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_d5eedfa744d4da30
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_d5eedfa744d4da30_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_0c22adf9c6a5bc0d.vhd when simulating
-- the core, cntr_11_0_0c22adf9c6a5bc0d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_0c22adf9c6a5bc0d IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END cntr_11_0_0c22adf9c6a5bc0d;

ARCHITECTURE cntr_11_0_0c22adf9c6a5bc0d_a OF cntr_11_0_0c22adf9c6a5bc0d IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_0c22adf9c6a5bc0d
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_0c22adf9c6a5bc0d USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 7,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_0c22adf9c6a5bc0d
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_0c22adf9c6a5bc0d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_6711bf92f3a48934.vhd when simulating
-- the core, bmg_72_6711bf92f3a48934. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_6711bf92f3a48934 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_6711bf92f3a48934;

ARCHITECTURE bmg_72_6711bf92f3a48934_a OF bmg_72_6711bf92f3a48934 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_6711bf92f3a48934
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_6711bf92f3a48934 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 7,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_6711bf92f3a48934.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 128,
      c_read_depth_b => 128,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 128,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_6711bf92f3a48934
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_6711bf92f3a48934_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_c8fdf7c1ceafa9d8.vhd when simulating
-- the core, addsb_11_0_c8fdf7c1ceafa9d8. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_c8fdf7c1ceafa9d8 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END addsb_11_0_c8fdf7c1ceafa9d8;

ARCHITECTURE addsb_11_0_c8fdf7c1ceafa9d8_a OF addsb_11_0_c8fdf7c1ceafa9d8 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_c8fdf7c1ceafa9d8
  PORT (
    a : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_c8fdf7c1ceafa9d8 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 3,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "000",
      c_b_width => 3,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 3,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_c8fdf7c1ceafa9d8
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_c8fdf7c1ceafa9d8_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_7e8fa68244af6cff.vhd when simulating
-- the core, bmg_72_7e8fa68244af6cff. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_7e8fa68244af6cff IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_7e8fa68244af6cff;

ARCHITECTURE bmg_72_7e8fa68244af6cff_a OF bmg_72_7e8fa68244af6cff IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_7e8fa68244af6cff
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_7e8fa68244af6cff USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 11,
      c_addrb_width => 11,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_7e8fa68244af6cff.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 2048,
      c_read_depth_b => 2048,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 2048,
      c_write_depth_b => 2048,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_7e8fa68244af6cff
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_7e8fa68244af6cff_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_1c323e86177437db.vhd when simulating
-- the core, dmg_72_1c323e86177437db. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_1c323e86177437db IS
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_1c323e86177437db;

ARCHITECTURE dmg_72_1c323e86177437db_a OF dmg_72_1c323e86177437db IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_1c323e86177437db
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_1c323e86177437db USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 5,
      c_default_data => "0",
      c_depth => 32,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_1c323e86177437db.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_1c323e86177437db
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_1c323e86177437db_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_070de696ab472038.vhd when simulating
-- the core, bmg_72_070de696ab472038. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_070de696ab472038 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_070de696ab472038;

ARCHITECTURE bmg_72_070de696ab472038_a OF bmg_72_070de696ab472038 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_070de696ab472038
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_070de696ab472038 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 8,
      c_addrb_width => 8,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_070de696ab472038.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 256,
      c_read_depth_b => 256,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 256,
      c_write_depth_b => 256,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_070de696ab472038
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_070de696ab472038_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_18f6f1cec46d694e.vhd when simulating
-- the core, addsb_11_0_18f6f1cec46d694e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_18f6f1cec46d694e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_18f6f1cec46d694e;

ARCHITECTURE addsb_11_0_18f6f1cec46d694e_a OF addsb_11_0_18f6f1cec46d694e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_18f6f1cec46d694e
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_18f6f1cec46d694e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_18f6f1cec46d694e
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_18f6f1cec46d694e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_ba1afd1a3b6d9138.vhd when simulating
-- the core, bmg_72_ba1afd1a3b6d9138. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_ba1afd1a3b6d9138 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_ba1afd1a3b6d9138;

ARCHITECTURE bmg_72_ba1afd1a3b6d9138_a OF bmg_72_ba1afd1a3b6d9138 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_ba1afd1a3b6d9138
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_ba1afd1a3b6d9138 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 5,
      c_addrb_width => 5,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_ba1afd1a3b6d9138.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 32,
      c_read_depth_b => 32,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 32,
      c_write_depth_b => 32,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_ba1afd1a3b6d9138
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_ba1afd1a3b6d9138_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_eb304381eda4ae1e.vhd when simulating
-- the core, bmg_72_eb304381eda4ae1e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_eb304381eda4ae1e IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_eb304381eda4ae1e;

ARCHITECTURE bmg_72_eb304381eda4ae1e_a OF bmg_72_eb304381eda4ae1e IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_eb304381eda4ae1e
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_eb304381eda4ae1e USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_eb304381eda4ae1e.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 64,
      c_read_depth_b => 64,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 64,
      c_write_depth_b => 64,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_eb304381eda4ae1e
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_eb304381eda4ae1e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_7789a80a5b2a8160.vhd when simulating
-- the core, cntr_11_0_7789a80a5b2a8160. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_7789a80a5b2a8160 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END cntr_11_0_7789a80a5b2a8160;

ARCHITECTURE cntr_11_0_7789a80a5b2a8160_a OF cntr_11_0_7789a80a5b2a8160 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_7789a80a5b2a8160
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_7789a80a5b2a8160 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 4,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_7789a80a5b2a8160
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_7789a80a5b2a8160_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_f0e087429b44571a.vhd when simulating
-- the core, bmg_72_f0e087429b44571a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_f0e087429b44571a IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_f0e087429b44571a;

ARCHITECTURE bmg_72_f0e087429b44571a_a OF bmg_72_f0e087429b44571a IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_f0e087429b44571a
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_f0e087429b44571a USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_f0e087429b44571a.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_f0e087429b44571a
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_f0e087429b44571a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_12b8e0a4a9ef4845.vhd when simulating
-- the core, cntr_11_0_12b8e0a4a9ef4845. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_12b8e0a4a9ef4845 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END cntr_11_0_12b8e0a4a9ef4845;

ARCHITECTURE cntr_11_0_12b8e0a4a9ef4845_a OF cntr_11_0_12b8e0a4a9ef4845 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_12b8e0a4a9ef4845
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_12b8e0a4a9ef4845 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_12b8e0a4a9ef4845
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_12b8e0a4a9ef4845_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_a1505185555f1882.vhd when simulating
-- the core, cntr_11_0_a1505185555f1882. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_a1505185555f1882 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END cntr_11_0_a1505185555f1882;

ARCHITECTURE cntr_11_0_a1505185555f1882_a OF cntr_11_0_a1505185555f1882 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_a1505185555f1882
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_a1505185555f1882 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 4,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_a1505185555f1882
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_a1505185555f1882_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_03f06ae367a98e8a.vhd when simulating
-- the core, cntr_11_0_03f06ae367a98e8a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_03f06ae367a98e8a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END cntr_11_0_03f06ae367a98e8a;

ARCHITECTURE cntr_11_0_03f06ae367a98e8a_a OF cntr_11_0_03f06ae367a98e8a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_03f06ae367a98e8a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_03f06ae367a98e8a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 7,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_03f06ae367a98e8a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_03f06ae367a98e8a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_4adf855dd0e5af2a.vhd when simulating
-- the core, cntr_11_0_4adf855dd0e5af2a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_4adf855dd0e5af2a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END cntr_11_0_4adf855dd0e5af2a;

ARCHITECTURE cntr_11_0_4adf855dd0e5af2a_a OF cntr_11_0_4adf855dd0e5af2a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_4adf855dd0e5af2a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_4adf855dd0e5af2a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 10,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_4adf855dd0e5af2a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_4adf855dd0e5af2a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_488bc588e4c66edf.vhd when simulating
-- the core, bmg_72_488bc588e4c66edf. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_488bc588e4c66edf IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_488bc588e4c66edf;

ARCHITECTURE bmg_72_488bc588e4c66edf_a OF bmg_72_488bc588e4c66edf IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_488bc588e4c66edf
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_488bc588e4c66edf USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 11,
      c_addrb_width => 11,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_488bc588e4c66edf.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 2048,
      c_read_depth_b => 2048,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 2048,
      c_write_depth_b => 2048,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_488bc588e4c66edf
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_488bc588e4c66edf_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_f54beabec7472b25.vhd when simulating
-- the core, dmg_72_f54beabec7472b25. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_f54beabec7472b25 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END dmg_72_f54beabec7472b25;

ARCHITECTURE dmg_72_f54beabec7472b25_a OF dmg_72_f54beabec7472b25 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_f54beabec7472b25
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_f54beabec7472b25 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 12,
      c_default_data => "0",
      c_depth => 4096,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_f54beabec7472b25.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 12
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_f54beabec7472b25
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_f54beabec7472b25_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_0b9daa5d24360c6e.vhd when simulating
-- the core, addsb_11_0_0b9daa5d24360c6e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_0b9daa5d24360c6e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_0b9daa5d24360c6e;

ARCHITECTURE addsb_11_0_0b9daa5d24360c6e_a OF addsb_11_0_0b9daa5d24360c6e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_0b9daa5d24360c6e
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_0b9daa5d24360c6e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_0b9daa5d24360c6e
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_0b9daa5d24360c6e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_d20b02a9f8239c7a.vhd when simulating
-- the core, dmg_72_d20b02a9f8239c7a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_d20b02a9f8239c7a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_d20b02a9f8239c7a;

ARCHITECTURE dmg_72_d20b02a9f8239c7a_a OF dmg_72_d20b02a9f8239c7a IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_d20b02a9f8239c7a
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_d20b02a9f8239c7a USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_d20b02a9f8239c7a.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_d20b02a9f8239c7a
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_d20b02a9f8239c7a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_533dcbdd307dbf50.vhd when simulating
-- the core, cntr_11_0_533dcbdd307dbf50. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_533dcbdd307dbf50 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END cntr_11_0_533dcbdd307dbf50;

ARCHITECTURE cntr_11_0_533dcbdd307dbf50_a OF cntr_11_0_533dcbdd307dbf50 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_533dcbdd307dbf50
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_533dcbdd307dbf50 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 2,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_533dcbdd307dbf50
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_533dcbdd307dbf50_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_60602034a1d84a16.vhd when simulating
-- the core, cntr_11_0_60602034a1d84a16. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_60602034a1d84a16 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
  );
END cntr_11_0_60602034a1d84a16;

ARCHITECTURE cntr_11_0_60602034a1d84a16_a OF cntr_11_0_60602034a1d84a16 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_60602034a1d84a16
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_60602034a1d84a16 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 11,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_60602034a1d84a16
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_60602034a1d84a16_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_b92ee532c1b215f1.vhd when simulating
-- the core, bmg_72_b92ee532c1b215f1. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_b92ee532c1b215f1 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_b92ee532c1b215f1;

ARCHITECTURE bmg_72_b92ee532c1b215f1_a OF bmg_72_b92ee532c1b215f1 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_b92ee532c1b215f1
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_b92ee532c1b215f1 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 7,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_b92ee532c1b215f1.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 128,
      c_read_depth_b => 128,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 128,
      c_write_depth_b => 128,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_b92ee532c1b215f1
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_b92ee532c1b215f1_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_505931c5b3ea228e.vhd when simulating
-- the core, dmg_72_505931c5b3ea228e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_505931c5b3ea228e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_505931c5b3ea228e;

ARCHITECTURE dmg_72_505931c5b3ea228e_a OF dmg_72_505931c5b3ea228e IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_505931c5b3ea228e
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_505931c5b3ea228e USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_505931c5b3ea228e.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_505931c5b3ea228e
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_505931c5b3ea228e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_9fff5a02c6b3c277.vhd when simulating
-- the core, bmg_72_9fff5a02c6b3c277. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_9fff5a02c6b3c277 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_9fff5a02c6b3c277;

ARCHITECTURE bmg_72_9fff5a02c6b3c277_a OF bmg_72_9fff5a02c6b3c277 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_9fff5a02c6b3c277
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_9fff5a02c6b3c277 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 9,
      c_addrb_width => 9,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_9fff5a02c6b3c277.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 512,
      c_read_depth_b => 512,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 512,
      c_write_depth_b => 512,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_9fff5a02c6b3c277
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_9fff5a02c6b3c277_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_b7550dc611e0410a.vhd when simulating
-- the core, cntr_11_0_b7550dc611e0410a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_b7550dc611e0410a IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_b7550dc611e0410a;

ARCHITECTURE cntr_11_0_b7550dc611e0410a_a OF cntr_11_0_b7550dc611e0410a IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_b7550dc611e0410a
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    load : IN STD_LOGIC;
    l : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_b7550dc611e0410a USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 1,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 1,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_b7550dc611e0410a
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    load => load,
    l => l,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_b7550dc611e0410a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_89850cbcf0fde6e9.vhd when simulating
-- the core, cntr_11_0_89850cbcf0fde6e9. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_89850cbcf0fde6e9 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END cntr_11_0_89850cbcf0fde6e9;

ARCHITECTURE cntr_11_0_89850cbcf0fde6e9_a OF cntr_11_0_89850cbcf0fde6e9 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_89850cbcf0fde6e9
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_89850cbcf0fde6e9 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 10,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_89850cbcf0fde6e9
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_89850cbcf0fde6e9_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_6bbb8fb0d8f20abe.vhd when simulating
-- the core, addsb_11_0_6bbb8fb0d8f20abe. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_6bbb8fb0d8f20abe IS
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END addsb_11_0_6bbb8fb0d8f20abe;

ARCHITECTURE addsb_11_0_6bbb8fb0d8f20abe_a OF addsb_11_0_6bbb8fb0d8f20abe IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_6bbb8fb0d8f20abe
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_6bbb8fb0d8f20abe USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 20,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000",
      c_b_width => 20,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 20,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_6bbb8fb0d8f20abe
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_6bbb8fb0d8f20abe_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_c9b173d075a3b6d7.vhd when simulating
-- the core, addsb_11_0_c9b173d075a3b6d7. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_c9b173d075a3b6d7 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_c9b173d075a3b6d7;

ARCHITECTURE addsb_11_0_c9b173d075a3b6d7_a OF addsb_11_0_c9b173d075a3b6d7 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_c9b173d075a3b6d7
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_c9b173d075a3b6d7 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_c9b173d075a3b6d7
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_c9b173d075a3b6d7_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_77dc1780892a0930.vhd when simulating
-- the core, bmg_72_77dc1780892a0930. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_77dc1780892a0930 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_77dc1780892a0930;

ARCHITECTURE bmg_72_77dc1780892a0930_a OF bmg_72_77dc1780892a0930 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_77dc1780892a0930
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_77dc1780892a0930 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_77dc1780892a0930.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_77dc1780892a0930
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_77dc1780892a0930_a;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
entity xlcounter_limit_fft_core is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned;
    cnt_63_48: integer:= 0;
    cnt_47_32: integer:= 0;
    cnt_31_16: integer:= 0;
    cnt_15_0: integer:= 0;
    count_limited: integer := 0
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_limit_fft_core ;
architecture behavior of xlcounter_limit_fft_core is
  signal high_cnt_to: std_logic_vector(31 downto 0);
  signal low_cnt_to: std_logic_vector(31 downto 0);
  signal cnt_to: std_logic_vector(63 downto 0);
  signal core_sinit, op_thresh0, core_ce: std_logic;
  signal rst_overrides_en: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
  -- synopsys translate_off
  signal real_op : real;
   -- synopsys translate_on
  function equals(op, cnt_to : std_logic_vector; width, arith : integer)
    return std_logic
  is
    variable signed_op, signed_cnt_to : signed (width - 1 downto 0);
    variable unsigned_op, unsigned_cnt_to : unsigned (width - 1 downto 0);
    variable result : std_logic;
  begin
    -- synopsys translate_off
    if ((is_XorU(op)) or (is_XorU(cnt_to)) ) then
      result := '0';
      return result;
    end if;
    -- synopsys translate_on
    if (op = cnt_to) then
      result := '1';
    else
      result := '0';
    end if;
    return result;
  end;
  component cntr_11_0_ed810b6704650710
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_ed810b6704650710:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_ed810b6704650710:
    component is "true";
  attribute box_type of cntr_11_0_ed810b6704650710:
    component  is "black_box";
  component cntr_11_0_125dc8e6a3ba8cad
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_125dc8e6a3ba8cad:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_125dc8e6a3ba8cad:
    component is "true";
  attribute box_type of cntr_11_0_125dc8e6a3ba8cad:
    component  is "black_box";
  component cntr_11_0_60602034a1d84a16
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_60602034a1d84a16:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_60602034a1d84a16:
    component is "true";
  attribute box_type of cntr_11_0_60602034a1d84a16:
    component  is "black_box";
  component cntr_11_0_89850cbcf0fde6e9
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_89850cbcf0fde6e9:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_89850cbcf0fde6e9:
    component is "true";
  attribute box_type of cntr_11_0_89850cbcf0fde6e9:
    component  is "black_box";
  component cntr_11_0_12b8e0a4a9ef4845
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_12b8e0a4a9ef4845:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_12b8e0a4a9ef4845:
    component is "true";
  attribute box_type of cntr_11_0_12b8e0a4a9ef4845:
    component  is "black_box";
  component cntr_11_0_133a8817831fb97a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_133a8817831fb97a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_133a8817831fb97a:
    component is "true";
  attribute box_type of cntr_11_0_133a8817831fb97a:
    component  is "black_box";
  component cntr_11_0_0c22adf9c6a5bc0d
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_0c22adf9c6a5bc0d:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_0c22adf9c6a5bc0d:
    component is "true";
  attribute box_type of cntr_11_0_0c22adf9c6a5bc0d:
    component  is "black_box";
  component cntr_11_0_d60ecc44fc05ecdd
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d60ecc44fc05ecdd:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d60ecc44fc05ecdd:
    component is "true";
  attribute box_type of cntr_11_0_d60ecc44fc05ecdd:
    component  is "black_box";
  component cntr_11_0_ee60311bb9d0db53
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_ee60311bb9d0db53:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_ee60311bb9d0db53:
    component is "true";
  attribute box_type of cntr_11_0_ee60311bb9d0db53:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec : std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec : std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
begin
  -- synopsys translate_off
  -- synopsys translate_on
  cnt_to(63 downto 48) <= integer_to_std_logic_vector(cnt_63_48, 16, op_arith);
  cnt_to(47 downto 32) <= integer_to_std_logic_vector(cnt_47_32, 16, op_arith);
  cnt_to(31 downto 16) <= integer_to_std_logic_vector(cnt_31_16, 16, op_arith);
  cnt_to(15 downto 0) <= integer_to_std_logic_vector(cnt_15_0, 16, op_arith);
  op <= op_net;
  core_ce <= ce and en(0);
  rst_overrides_en <= rst(0) or en(0);
  limit : if (count_limited = 1) generate
    eq_cnt_to : process (op_net, cnt_to)
    begin
      op_thresh0 <= equals(op_net, cnt_to(op_width - 1 downto 0),
                     op_width, op_arith);
    end process;
    core_sinit <= (op_thresh0 or clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  no_limit : if (count_limited = 0) generate
    core_sinit <= (clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  comp0: if ((core_name0 = "cntr_11_0_ed810b6704650710")) generate
    core_instance0: cntr_11_0_ed810b6704650710
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_125dc8e6a3ba8cad")) generate
    core_instance1: cntr_11_0_125dc8e6a3ba8cad
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp2: if ((core_name0 = "cntr_11_0_60602034a1d84a16")) generate
    core_instance2: cntr_11_0_60602034a1d84a16
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp3: if ((core_name0 = "cntr_11_0_89850cbcf0fde6e9")) generate
    core_instance3: cntr_11_0_89850cbcf0fde6e9
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp4: if ((core_name0 = "cntr_11_0_12b8e0a4a9ef4845")) generate
    core_instance4: cntr_11_0_12b8e0a4a9ef4845
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp5: if ((core_name0 = "cntr_11_0_133a8817831fb97a")) generate
    core_instance5: cntr_11_0_133a8817831fb97a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp6: if ((core_name0 = "cntr_11_0_0c22adf9c6a5bc0d")) generate
    core_instance6: cntr_11_0_0c22adf9c6a5bc0d
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp7: if ((core_name0 = "cntr_11_0_d60ecc44fc05ecdd")) generate
    core_instance7: cntr_11_0_d60ecc44fc05ecdd
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp8: if ((core_name0 = "cntr_11_0_ee60311bb9d0db53")) generate
    core_instance8: cntr_11_0_ee60311bb9d0db53
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlspram_fft_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
    );
  port (
    data_in: in std_logic_vector(c_width - 1 downto 0);
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    we: in std_logic_vector(0 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data_out: out std_logic_vector(c_width - 1 downto 0)
  );
end xlspram_fft_core ;
architecture behavior of xlspram_fft_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_data_out, dly_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_we, core_ce, sinit: std_logic;
  component bmg_72_77dc1780892a0930
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_77dc1780892a0930:
    component is true;
  attribute fpga_dont_touch of bmg_72_77dc1780892a0930:
    component is "true";
  attribute box_type of bmg_72_77dc1780892a0930:
    component  is "black_box";
  component bmg_72_f0e087429b44571a
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_f0e087429b44571a:
    component is true;
  attribute fpga_dont_touch of bmg_72_f0e087429b44571a:
    component is "true";
  attribute box_type of bmg_72_f0e087429b44571a:
    component  is "black_box";
  component bmg_72_7e8fa68244af6cff
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_7e8fa68244af6cff:
    component is true;
  attribute fpga_dont_touch of bmg_72_7e8fa68244af6cff:
    component is "true";
  attribute box_type of bmg_72_7e8fa68244af6cff:
    component  is "black_box";
  component bmg_72_756e5f183b33a31a
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_756e5f183b33a31a:
    component is true;
  attribute fpga_dont_touch of bmg_72_756e5f183b33a31a:
    component is "true";
  attribute box_type of bmg_72_756e5f183b33a31a:
    component  is "black_box";
  component bmg_72_9fff5a02c6b3c277
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_9fff5a02c6b3c277:
    component is true;
  attribute fpga_dont_touch of bmg_72_9fff5a02c6b3c277:
    component is "true";
  attribute box_type of bmg_72_9fff5a02c6b3c277:
    component  is "black_box";
  component bmg_72_87bb354a843dab37
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_87bb354a843dab37:
    component is true;
  attribute fpga_dont_touch of bmg_72_87bb354a843dab37:
    component is "true";
  attribute box_type of bmg_72_87bb354a843dab37:
    component  is "black_box";
  component bmg_72_b92ee532c1b215f1
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_b92ee532c1b215f1:
    component is true;
  attribute fpga_dont_touch of bmg_72_b92ee532c1b215f1:
    component is "true";
  attribute box_type of bmg_72_b92ee532c1b215f1:
    component  is "black_box";
  component bmg_72_59143b4ed22b761d
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_59143b4ed22b761d:
    component is true;
  attribute fpga_dont_touch of bmg_72_59143b4ed22b761d:
    component is "true";
  attribute box_type of bmg_72_59143b4ed22b761d:
    component  is "black_box";
  component bmg_72_ba1afd1a3b6d9138
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_ba1afd1a3b6d9138:
    component is true;
  attribute fpga_dont_touch of bmg_72_ba1afd1a3b6d9138:
    component is "true";
  attribute box_type of bmg_72_ba1afd1a3b6d9138:
    component  is "black_box";
begin
  data_out <= dly_data_out;
  core_we <= we(0);
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_77dc1780892a0930")) generate
    core_instance0: bmg_72_77dc1780892a0930
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_f0e087429b44571a")) generate
    core_instance1: bmg_72_f0e087429b44571a
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp2: if ((core_name0 = "bmg_72_7e8fa68244af6cff")) generate
    core_instance2: bmg_72_7e8fa68244af6cff
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp3: if ((core_name0 = "bmg_72_756e5f183b33a31a")) generate
    core_instance3: bmg_72_756e5f183b33a31a
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp4: if ((core_name0 = "bmg_72_9fff5a02c6b3c277")) generate
    core_instance4: bmg_72_9fff5a02c6b3c277
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp5: if ((core_name0 = "bmg_72_87bb354a843dab37")) generate
    core_instance5: bmg_72_87bb354a843dab37
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp6: if ((core_name0 = "bmg_72_b92ee532c1b215f1")) generate
    core_instance6: bmg_72_b92ee532c1b215f1
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp7: if ((core_name0 = "bmg_72_59143b4ed22b761d")) generate
    core_instance7: bmg_72_59143b4ed22b761d
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp8: if ((core_name0 = "bmg_72_ba1afd1a3b6d9138")) generate
    core_instance8: bmg_72_ba1afd1a3b6d9138
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => dly_data_out
      );
  end generate;
  latency_1: if (latency <= 1) generate
    dly_data_out <= core_data_out;
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9a0fa0f632 is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9a0fa0f632;


architecture behavior of reinterpret_9a0fa0f632 is
  signal input_port_1_40: unsigned((18 - 1) downto 0);
  signal output_port_5_5_force: signed((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlslice is
    generic (
        new_msb      : integer := 9;
        new_lsb      : integer := 1;
        x_width      : integer := 16;
        y_width      : integer := 8);
    port (
        x : in std_logic_vector (x_width-1 downto 0);
        y : out std_logic_vector (y_width-1 downto 0));
end xlslice;
architecture behavior of xlslice is
begin
    y <= x(new_msb downto new_lsb);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_bc4405cd1e is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_bc4405cd1e;


architecture behavior of reinterpret_bc4405cd1e is
  signal input_port_1_40: signed((19 - 1) downto 0);
  signal output_port_5_5_force: unsigned((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub_fft_core is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub_fft_core;
architecture behavior of xladdsub_fft_core is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_59920783799a8e86
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_18f6f1cec46d694e
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_0b9daa5d24360c6e
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_c9b173d075a3b6d7
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_6bbb8fb0d8f20abe
    port (
          a: in std_logic_vector(20 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(20 - 1 downto 0)
    );
  end component;
  component addsb_11_0_a0497faccc62b6b2
    port (
          a: in std_logic_vector(20 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(20 - 1 downto 0)
    );
  end component;
  component addsb_11_0_c8fdf7c1ceafa9d8
    port (
          a: in std_logic_vector(3 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(3 - 1 downto 0)
    );
  end component;
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_59920783799a8e86")) generate
    core_instance0: addsb_11_0_59920783799a8e86
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp1: if ((core_name0 = "addsb_11_0_18f6f1cec46d694e")) generate
    core_instance1: addsb_11_0_18f6f1cec46d694e
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_0b9daa5d24360c6e")) generate
    core_instance2: addsb_11_0_0b9daa5d24360c6e
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp3: if ((core_name0 = "addsb_11_0_c9b173d075a3b6d7")) generate
    core_instance3: addsb_11_0_c9b173d075a3b6d7
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp4: if ((core_name0 = "addsb_11_0_6bbb8fb0d8f20abe")) generate
    core_instance4: addsb_11_0_6bbb8fb0d8f20abe
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp5: if ((core_name0 = "addsb_11_0_a0497faccc62b6b2")) generate
    core_instance5: addsb_11_0_a0497faccc62b6b2
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp6: if ((core_name0 = "addsb_11_0_c8fdf7c1ceafa9d8")) generate
    core_instance6: addsb_11_0_c8fdf7c1ceafa9d8
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a246e373e7 is
  port (
    in0 : in std_logic_vector((18 - 1) downto 0);
    in1 : in std_logic_vector((18 - 1) downto 0);
    in2 : in std_logic_vector((18 - 1) downto 0);
    in3 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((72 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a246e373e7;


architecture behavior of concat_a246e373e7 is
  signal in0_1_23: unsigned((18 - 1) downto 0);
  signal in1_1_27: unsigned((18 - 1) downto 0);
  signal in2_1_31: unsigned((18 - 1) downto 0);
  signal in3_1_35: unsigned((18 - 1) downto 0);
  signal y_2_1_concat: unsigned((72 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_580feec131 is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_580feec131;


architecture behavior of reinterpret_580feec131 is
  signal input_port_1_40: signed((18 - 1) downto 0);
  signal output_port_5_5_force: unsigned((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_504cae28bd is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_504cae28bd;


architecture behavior of concat_504cae28bd is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((20 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_f4186754a0 is
  port (
    a : in std_logic_vector((20 - 1) downto 0);
    b : in std_logic_vector((19 - 1) downto 0);
    s : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_f4186754a0;


architecture behavior of addsub_f4186754a0 is
  signal a_17_32: signed((20 - 1) downto 0);
  signal b_17_35: unsigned((19 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (3 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_91_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_91_20_back: signed((18 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (3 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((21 - 1) downto 0);
  signal cast_69_22: signed((21 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((21 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((18 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(2);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(2);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 2 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 19, 21, 19);
  cast_69_22 <= u2s_cast(b_17_35, 19, 21, 19);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 19, 18, 17);
  op_mem_91_20_front_din <= cast_internal_s_83_3_convert;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4709ea49b5 is
  port (
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4709ea49b5;


architecture behavior of constant_4709ea49b5 is
begin
  op <= "0000000000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_f661f8d9b7 is
  port (
    input_port : in std_logic_vector((20 - 1) downto 0);
    output_port : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_f661f8d9b7;


architecture behavior of reinterpret_f661f8d9b7 is
  signal input_port_1_40: unsigned((20 - 1) downto 0);
  signal output_port_5_5_force: signed((20 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d2180c9169 is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d2180c9169;


architecture behavior of reinterpret_d2180c9169 is
  signal input_port_1_40: unsigned((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_938d99ac11 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_938d99ac11;


architecture behavior of logical_938d99ac11 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_63700884f5 is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_63700884f5;


architecture behavior of reinterpret_63700884f5 is
  signal input_port_1_40: unsigned((19 - 1) downto 0);
  signal output_port_5_5_force: signed((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9306b5127f is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9306b5127f;


architecture behavior of reinterpret_9306b5127f is
  signal input_port_1_40: unsigned((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2aea51ccde is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((19 - 1) downto 0);
    in2 : in std_logic_vector((19 - 1) downto 0);
    in3 : in std_logic_vector((19 - 1) downto 0);
    y : out std_logic_vector((76 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2aea51ccde;


architecture behavior of concat_2aea51ccde is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((19 - 1) downto 0);
  signal in2_1_31: unsigned((19 - 1) downto 0);
  signal in3_1_35: unsigned((19 - 1) downto 0);
  signal y_2_1_concat: unsigned((76 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity scale_9f61027ba4 is
  port (
    ip : in std_logic_vector((19 - 1) downto 0);
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end scale_9f61027ba4;


architecture behavior of scale_9f61027ba4 is
  signal ip_17_23: signed((19 - 1) downto 0);
begin
  ip_17_23 <= std_logic_vector_to_signed(ip);
  op <= signed_to_std_logic_vector(ip_17_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_b198bd62b0 is
  port (
    in0 : in std_logic_vector((18 - 1) downto 0);
    in1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_b198bd62b0;


architecture behavior of concat_b198bd62b0 is
  signal in0_1_23: unsigned((18 - 1) downto 0);
  signal in1_1_27: unsigned((18 - 1) downto 0);
  signal y_2_1_concat: unsigned((36 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_86b044698f is
  port (
    input_port : in std_logic_vector((36 - 1) downto 0);
    output_port : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_86b044698f;


architecture behavior of reinterpret_86b044698f is
  signal input_port_1_40: unsigned((36 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_f983e30a8b is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_f983e30a8b;


architecture behavior of negate_f983e30a8b is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (1 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    0 => "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal cast_internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(0);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  cast_internal_ip_40_3_convert <= s2s_cast(internal_ip_join_30_1, 17, 18, 17);
  op_mem_48_20_push_front_pop_back_en <= '0';
  op <= signed_to_std_logic_vector(cast_internal_ip_40_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_6699ee0916 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_6699ee0916;


architecture behavior of delay_6699ee0916 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e47f8076b8 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e47f8076b8;


architecture behavior of constant_e47f8076b8 is
begin
  op <= "1000000000000";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlcounter_free_fft_core is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free_fft_core ;
architecture behavior of xlcounter_free_fft_core is
  component cntr_11_0_125dc8e6a3ba8cad
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_125dc8e6a3ba8cad:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_125dc8e6a3ba8cad:
    component is "true";
  attribute box_type of cntr_11_0_125dc8e6a3ba8cad:
    component  is "black_box";
  component cntr_11_0_461fd5d45cff2f9b
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_461fd5d45cff2f9b:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_461fd5d45cff2f9b:
    component is "true";
  attribute box_type of cntr_11_0_461fd5d45cff2f9b:
    component  is "black_box";
  component cntr_11_0_ed810b6704650710
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_ed810b6704650710:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_ed810b6704650710:
    component is "true";
  attribute box_type of cntr_11_0_ed810b6704650710:
    component  is "black_box";
  component cntr_11_0_a1505185555f1882
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_a1505185555f1882:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_a1505185555f1882:
    component is "true";
  attribute box_type of cntr_11_0_a1505185555f1882:
    component  is "black_box";
  component cntr_11_0_7789a80a5b2a8160
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_7789a80a5b2a8160:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_7789a80a5b2a8160:
    component is "true";
  attribute box_type of cntr_11_0_7789a80a5b2a8160:
    component  is "black_box";
  component cntr_11_0_3a3ea2f70b8548a5
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_3a3ea2f70b8548a5:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_3a3ea2f70b8548a5:
    component is "true";
  attribute box_type of cntr_11_0_3a3ea2f70b8548a5:
    component  is "black_box";
  component cntr_11_0_efa60dbe2ed9d35a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_efa60dbe2ed9d35a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_efa60dbe2ed9d35a:
    component is "true";
  attribute box_type of cntr_11_0_efa60dbe2ed9d35a:
    component  is "black_box";
  component cntr_11_0_99383d874600f8be
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_99383d874600f8be:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_99383d874600f8be:
    component is "true";
  attribute box_type of cntr_11_0_99383d874600f8be:
    component  is "black_box";
  component cntr_11_0_533dcbdd307dbf50
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_533dcbdd307dbf50:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_533dcbdd307dbf50:
    component is "true";
  attribute box_type of cntr_11_0_533dcbdd307dbf50:
    component  is "black_box";
  component cntr_11_0_a2916e7e77833dd6
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_a2916e7e77833dd6:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_a2916e7e77833dd6:
    component is "true";
  attribute box_type of cntr_11_0_a2916e7e77833dd6:
    component  is "black_box";
  component cntr_11_0_2f7113c203379501
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_2f7113c203379501:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_2f7113c203379501:
    component is "true";
  attribute box_type of cntr_11_0_2f7113c203379501:
    component  is "black_box";
  component cntr_11_0_60602034a1d84a16
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_60602034a1d84a16:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_60602034a1d84a16:
    component is "true";
  attribute box_type of cntr_11_0_60602034a1d84a16:
    component  is "black_box";
  component cntr_11_0_4adf855dd0e5af2a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_4adf855dd0e5af2a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_4adf855dd0e5af2a:
    component is "true";
  attribute box_type of cntr_11_0_4adf855dd0e5af2a:
    component  is "black_box";
  component cntr_11_0_89850cbcf0fde6e9
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_89850cbcf0fde6e9:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_89850cbcf0fde6e9:
    component is "true";
  attribute box_type of cntr_11_0_89850cbcf0fde6e9:
    component  is "black_box";
  component cntr_11_0_796a9d3dfbc0c498
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_796a9d3dfbc0c498:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_796a9d3dfbc0c498:
    component is "true";
  attribute box_type of cntr_11_0_796a9d3dfbc0c498:
    component  is "black_box";
  component cntr_11_0_12b8e0a4a9ef4845
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_12b8e0a4a9ef4845:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_12b8e0a4a9ef4845:
    component is "true";
  attribute box_type of cntr_11_0_12b8e0a4a9ef4845:
    component  is "black_box";
  component cntr_11_0_b7550dc611e0410a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_b7550dc611e0410a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_b7550dc611e0410a:
    component is "true";
  attribute box_type of cntr_11_0_b7550dc611e0410a:
    component  is "black_box";
  component cntr_11_0_133a8817831fb97a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_133a8817831fb97a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_133a8817831fb97a:
    component is "true";
  attribute box_type of cntr_11_0_133a8817831fb97a:
    component  is "black_box";
  component cntr_11_0_03f06ae367a98e8a
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_03f06ae367a98e8a:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_03f06ae367a98e8a:
    component is "true";
  attribute box_type of cntr_11_0_03f06ae367a98e8a:
    component  is "black_box";
  component cntr_11_0_0c22adf9c6a5bc0d
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_0c22adf9c6a5bc0d:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_0c22adf9c6a5bc0d:
    component is "true";
  attribute box_type of cntr_11_0_0c22adf9c6a5bc0d:
    component  is "black_box";
  component cntr_11_0_cb1ffe90ceffe54f
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_cb1ffe90ceffe54f:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_cb1ffe90ceffe54f:
    component is "true";
  attribute box_type of cntr_11_0_cb1ffe90ceffe54f:
    component  is "black_box";
  component cntr_11_0_d60ecc44fc05ecdd
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d60ecc44fc05ecdd:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d60ecc44fc05ecdd:
    component is "true";
  attribute box_type of cntr_11_0_d60ecc44fc05ecdd:
    component  is "black_box";
  component cntr_11_0_d5eedfa744d4da30
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      load: in std_logic;
      l: in std_logic_vector(op_width - 1 downto 0);
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d5eedfa744d4da30:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d5eedfa744d4da30:
    component is "true";
  attribute box_type of cntr_11_0_d5eedfa744d4da30:
    component  is "black_box";
  component cntr_11_0_ee60311bb9d0db53
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_ee60311bb9d0db53:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_ee60311bb9d0db53:
    component is "true";
  attribute box_type of cntr_11_0_ee60311bb9d0db53:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_125dc8e6a3ba8cad")) generate
    core_instance0: cntr_11_0_125dc8e6a3ba8cad
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_461fd5d45cff2f9b")) generate
    core_instance1: cntr_11_0_461fd5d45cff2f9b
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp2: if ((core_name0 = "cntr_11_0_ed810b6704650710")) generate
    core_instance2: cntr_11_0_ed810b6704650710
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp3: if ((core_name0 = "cntr_11_0_a1505185555f1882")) generate
    core_instance3: cntr_11_0_a1505185555f1882
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp4: if ((core_name0 = "cntr_11_0_7789a80a5b2a8160")) generate
    core_instance4: cntr_11_0_7789a80a5b2a8160
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp5: if ((core_name0 = "cntr_11_0_3a3ea2f70b8548a5")) generate
    core_instance5: cntr_11_0_3a3ea2f70b8548a5
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp6: if ((core_name0 = "cntr_11_0_efa60dbe2ed9d35a")) generate
    core_instance6: cntr_11_0_efa60dbe2ed9d35a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp7: if ((core_name0 = "cntr_11_0_99383d874600f8be")) generate
    core_instance7: cntr_11_0_99383d874600f8be
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp8: if ((core_name0 = "cntr_11_0_533dcbdd307dbf50")) generate
    core_instance8: cntr_11_0_533dcbdd307dbf50
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp9: if ((core_name0 = "cntr_11_0_a2916e7e77833dd6")) generate
    core_instance9: cntr_11_0_a2916e7e77833dd6
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp10: if ((core_name0 = "cntr_11_0_2f7113c203379501")) generate
    core_instance10: cntr_11_0_2f7113c203379501
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp11: if ((core_name0 = "cntr_11_0_60602034a1d84a16")) generate
    core_instance11: cntr_11_0_60602034a1d84a16
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp12: if ((core_name0 = "cntr_11_0_4adf855dd0e5af2a")) generate
    core_instance12: cntr_11_0_4adf855dd0e5af2a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp13: if ((core_name0 = "cntr_11_0_89850cbcf0fde6e9")) generate
    core_instance13: cntr_11_0_89850cbcf0fde6e9
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp14: if ((core_name0 = "cntr_11_0_796a9d3dfbc0c498")) generate
    core_instance14: cntr_11_0_796a9d3dfbc0c498
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp15: if ((core_name0 = "cntr_11_0_12b8e0a4a9ef4845")) generate
    core_instance15: cntr_11_0_12b8e0a4a9ef4845
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp16: if ((core_name0 = "cntr_11_0_b7550dc611e0410a")) generate
    core_instance16: cntr_11_0_b7550dc611e0410a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp17: if ((core_name0 = "cntr_11_0_133a8817831fb97a")) generate
    core_instance17: cntr_11_0_133a8817831fb97a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp18: if ((core_name0 = "cntr_11_0_03f06ae367a98e8a")) generate
    core_instance18: cntr_11_0_03f06ae367a98e8a
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp19: if ((core_name0 = "cntr_11_0_0c22adf9c6a5bc0d")) generate
    core_instance19: cntr_11_0_0c22adf9c6a5bc0d
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp20: if ((core_name0 = "cntr_11_0_cb1ffe90ceffe54f")) generate
    core_instance20: cntr_11_0_cb1ffe90ceffe54f
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp21: if ((core_name0 = "cntr_11_0_d60ecc44fc05ecdd")) generate
    core_instance21: cntr_11_0_d60ecc44fc05ecdd
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp22: if ((core_name0 = "cntr_11_0_d5eedfa744d4da30")) generate
    core_instance22: cntr_11_0_d5eedfa744d4da30
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        load => load(0),
        l => din,
        q => op_net
      );
  end generate;
  comp23: if ((core_name0 = "cntr_11_0_ee60311bb9d0db53")) generate
    core_instance23: cntr_11_0_ee60311bb9d0db53
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_bdaf6c9e55 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_bdaf6c9e55;


architecture behavior of delay_bdaf6c9e55 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (4 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(3);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_fca786f2ff is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((36 - 1) downto 0);
    d1 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_fca786f2ff;


architecture behavior of mux_fca786f2ff is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((36 - 1) downto 0);
  signal d1_1_27: std_logic_vector((36 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((36 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_54e7975215 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54e7975215;


architecture behavior of relational_54e7975215 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_c53de546ea is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_c53de546ea;


architecture behavior of delay_c53de546ea is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (4 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(3);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_9f02caa990 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_9f02caa990;


architecture behavior of delay_9f02caa990 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_50be3b5040 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_50be3b5040;


architecture behavior of constant_50be3b5040 is
begin
  op <= "0000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0c8736a503 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0c8736a503;


architecture behavior of constant_0c8736a503 is
begin
  op <= "0000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_80f90b97d0 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_80f90b97d0;


architecture behavior of logical_80f90b97d0 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1bef4ba0e4 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1bef4ba0e4;


architecture behavior of mux_1bef4ba0e4 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal unregy_join_6_1: std_logic;
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= std_logic_to_vector(unregy_join_6_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6dfa374756 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6dfa374756;


architecture behavior of relational_6dfa374756 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2550da35d2 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2550da35d2;


architecture behavior of relational_2550da35d2 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_25f2d74a2a is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_25f2d74a2a;


architecture behavior of mux_25f2d74a2a is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000");
  signal pipe_16_22_front_din: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4670f4967f is
  port (
    d : in std_logic_vector((12 - 1) downto 0);
    q : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4670f4967f;


architecture behavior of delay_4670f4967f is
  signal d_1_22: std_logic_vector((12 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e4b9fcaf02 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e4b9fcaf02;


architecture behavior of delay_e4b9fcaf02 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_21355083c1 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_21355083c1;


architecture behavior of delay_21355083c1 is
  signal d_1_22: std_logic_vector((1 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_dist_fft_core is
  generic (
    core_name0: string := "";
    addr_width: integer := 2;
    latency: integer := 0;
    c_width: integer := 12;
    c_address_width: integer := 4
  );
  port (
    addr: in std_logic_vector(addr_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_dist_fft_core ;
architecture behavior of xlsprom_dist_fft_core is
  component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i           : in std_logic_vector(width - 1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width - 1 downto 0));
  end component;
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  constant num_extra_addr_bits: integer := (c_address_width - addr_width);
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_ce: std_logic;
  component dmg_72_08915946f5ebdf9c
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_08915946f5ebdf9c:
    component is true;
  attribute fpga_dont_touch of dmg_72_08915946f5ebdf9c:
    component is "true";
  attribute box_type of dmg_72_08915946f5ebdf9c:
    component  is "black_box";
  component dmg_72_b5cea772b1c370b5
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_b5cea772b1c370b5:
    component is true;
  attribute fpga_dont_touch of dmg_72_b5cea772b1c370b5:
    component is "true";
  attribute box_type of dmg_72_b5cea772b1c370b5:
    component  is "black_box";
  component dmg_72_f54beabec7472b25
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_f54beabec7472b25:
    component is true;
  attribute fpga_dont_touch of dmg_72_f54beabec7472b25:
    component is "true";
  attribute box_type of dmg_72_f54beabec7472b25:
    component  is "black_box";
begin
  need_to_pad_addr: if num_extra_addr_bits > 0 generate
      core_addr(c_address_width - 1 downto addr_width) <= (others => '0');
    core_addr(addr_width - 1 downto 0) <= addr;
  end generate;
  no_need_to_pad_addr: if num_extra_addr_bits = 0 generate
    core_addr <= addr;
  end generate;
  core_ce <= ce and en(0);
  comp0: if ((core_name0 = "dmg_72_08915946f5ebdf9c")) generate
    core_instance0: dmg_72_08915946f5ebdf9c
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp1: if ((core_name0 = "dmg_72_b5cea772b1c370b5")) generate
    core_instance1: dmg_72_b5cea772b1c370b5
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp2: if ((core_name0 = "dmg_72_f54beabec7472b25")) generate
    core_instance2: dmg_72_f54beabec7472b25
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_0_or_1: if (latency <= 1)
  generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_23d71a76f2 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_23d71a76f2;


architecture behavior of delay_23d71a76f2 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_aab7b18c27 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_aab7b18c27;


architecture behavior of delay_aab7b18c27 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (6 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(5);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_5a12f8f9be is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((19 - 1) downto 0);
    y : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_5a12f8f9be;


architecture behavior of concat_5a12f8f9be is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((19 - 1) downto 0);
  signal y_2_1_concat: unsigned((38 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c615d93998 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c615d93998;


architecture behavior of concat_c615d93998 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((21 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_4a8cbc85ce is
  port (
    input_port : in std_logic_vector((20 - 1) downto 0);
    output_port : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_4a8cbc85ce;


architecture behavior of reinterpret_4a8cbc85ce is
  signal input_port_1_40: signed((20 - 1) downto 0);
  signal output_port_5_5_force: unsigned((20 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_b96bfee539 is
  port (
    a : in std_logic_vector((21 - 1) downto 0);
    b : in std_logic_vector((19 - 1) downto 0);
    s : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_b96bfee539;


architecture behavior of addsub_b96bfee539 is
  signal a_17_32: signed((21 - 1) downto 0);
  signal b_17_35: unsigned((19 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (3 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_91_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_91_20_back: signed((18 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (3 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((22 - 1) downto 0);
  signal cast_69_22: signed((22 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((22 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((18 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(2);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(2);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 2 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 19, 22, 19);
  cast_69_22 <= u2s_cast(b_17_35, 19, 22, 19);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 19, 18, 17);
  op_mem_91_20_front_din <= cast_internal_s_83_3_convert;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d357e69fa3 is
  port (
    input_port : in std_logic_vector((21 - 1) downto 0);
    output_port : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d357e69fa3;


architecture behavior of reinterpret_d357e69fa3 is
  signal input_port_1_40: unsigned((21 - 1) downto 0);
  signal output_port_5_5_force: signed((21 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_9d76333483 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_9d76333483;


architecture behavior of logical_9d76333483 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_5bc1b3bb27 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_5bc1b3bb27;


architecture behavior of logical_5bc1b3bb27 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (3 - 1)) of std_logic;
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    '0',
    '0',
    '0');
  signal latency_pipe_5_26_front_din: std_logic;
  signal latency_pipe_5_26_back: std_logic;
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal bit_2_27: std_logic;
  signal fully_2_1_bitnot: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(2);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          latency_pipe_5_26(i) <= latency_pipe_5_26(i-1);
        end loop;
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  bit_2_27 <= d0_1_24 and d1_1_27;
  fully_2_1_bitnot <= not bit_2_27;
  latency_pipe_5_26_front_din <= fully_2_1_bitnot;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= std_logic_to_vector(latency_pipe_5_26_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0c7cd7a34 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0c7cd7a34;


architecture behavior of concat_a0c7cd7a34 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_112d91c147 is
  port (
    input_port : in std_logic_vector((1 - 1) downto 0);
    output_port : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_112d91c147;


architecture behavior of reinterpret_112d91c147 is
  signal input_port_1_40: boolean;
  signal output_port_7_5_convert: unsigned((1 - 1) downto 0);
begin
  input_port_1_40 <= ((input_port) = "1");
  output_port_7_5_convert <= u2u_cast(std_logic_vector_to_unsigned(boolean_to_vector(input_port_1_40)), 0, 1, 0);
  output_port <= unsigned_to_std_logic_vector(output_port_7_5_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_f86ebb6084 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((20 - 1) downto 0);
    in2 : in std_logic_vector((20 - 1) downto 0);
    in3 : in std_logic_vector((20 - 1) downto 0);
    y : out std_logic_vector((80 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_f86ebb6084;


architecture behavior of concat_f86ebb6084 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((20 - 1) downto 0);
  signal in2_1_31: unsigned((20 - 1) downto 0);
  signal in3_1_35: unsigned((20 - 1) downto 0);
  signal y_2_1_concat: unsigned((80 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_ba2df6ec2d is
  port (
    a : in std_logic_vector((20 - 1) downto 0);
    b : in std_logic_vector((19 - 1) downto 0);
    s : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_ba2df6ec2d;


architecture behavior of addsub_ba2df6ec2d is
  signal a_17_32: signed((20 - 1) downto 0);
  signal b_17_35: unsigned((19 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (1 - 1)) of signed((20 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    0 => "00000000000000000000");
  signal op_mem_91_20_front_din: signed((20 - 1) downto 0);
  signal op_mem_91_20_back: signed((20 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (1 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    0 => "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((21 - 1) downto 0);
  signal cast_69_22: signed((21 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((21 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((20 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(0);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(0);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 19, 21, 19);
  cast_69_22 <= u2s_cast(b_17_35, 19, 21, 19);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 19, 20, 18);
  op_mem_91_20_push_front_pop_back_en <= '0';
  cout_mem_92_22_push_front_pop_back_en <= '0';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(cast_internal_s_83_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b366689086 is
  port (
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b366689086;


architecture behavior of constant_b366689086 is
begin
  op <= "0000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_b1e9d7c303 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_b1e9d7c303;


architecture behavior of logical_b1e9d7c303 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal bit_2_26: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bitnot: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  bit_2_26 <= d0_1_24 or d1_1_27;
  fully_2_1_bitnot <= not bit_2_26;
  y <= fully_2_1_bitnot;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d610556e85 is
  port (
    input_port : in std_logic_vector((4 - 1) downto 0);
    output_port : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d610556e85;


architecture behavior of reinterpret_d610556e85 is
  signal input_port_1_40: unsigned((4 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_d930162434 is
  port (
    a : in std_logic_vector((4 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_d930162434;


architecture behavior of relational_d930162434 is
  signal a_1_31: unsigned((4 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_bd20dd351d is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_bd20dd351d;


architecture behavior of concat_bd20dd351d is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((2 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9a54e08c7c is
  port (
    input_port : in std_logic_vector((2 - 1) downto 0);
    output_port : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9a54e08c7c;


architecture behavior of reinterpret_9a54e08c7c is
  signal input_port_1_40: unsigned((2 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4822199898 is
  port (
    in0 : in std_logic_vector((38 - 1) downto 0);
    in1 : in std_logic_vector((38 - 1) downto 0);
    y : out std_logic_vector((76 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4822199898;


architecture behavior of concat_4822199898 is
  signal in0_1_23: unsigned((38 - 1) downto 0);
  signal in1_1_27: unsigned((38 - 1) downto 0);
  signal y_2_1_concat: unsigned((76 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_9ff8aec2dc is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((80 - 1) downto 0);
    d1 : in std_logic_vector((80 - 1) downto 0);
    y : out std_logic_vector((80 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_9ff8aec2dc;


architecture behavior of mux_9ff8aec2dc is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((80 - 1) downto 0);
  signal d1_1_27: std_logic_vector((80 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((80 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((80 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((80 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((80 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4c449dd556 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4c449dd556;


architecture behavior of constant_4c449dd556 is
begin
  op <= "0000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_fa260f7d22 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_fa260f7d22;


architecture behavior of delay_fa260f7d22 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (7 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(6);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 6 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e18fb31a3d is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e18fb31a3d;


architecture behavior of delay_e18fb31a3d is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_0309b30f97 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_0309b30f97;


architecture behavior of logical_0309b30f97 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  type array_type_latency_pipe_5_26 is array (0 to (1 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    0 => "0");
  signal latency_pipe_5_26_front_din: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_back: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  latency_pipe_5_26_back <= latency_pipe_5_26(0);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  latency_pipe_5_26_front_din <= fully_2_1_bit;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= latency_pipe_5_26_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4bb6f691f7 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((36 - 1) downto 0);
    d1 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4bb6f691f7;


architecture behavior of mux_4bb6f691f7 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((36 - 1) downto 0);
  signal d1_1_27: std_logic_vector((36 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((36 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9e724c4b50 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((20 - 1) downto 0);
    y : out std_logic_vector((40 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9e724c4b50;


architecture behavior of concat_9e724c4b50 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((20 - 1) downto 0);
  signal y_2_1_concat: unsigned((40 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e6bc20c81b is
  port (
    in0 : in std_logic_vector((21 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((22 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e6bc20c81b;


architecture behavior of concat_e6bc20c81b is
  signal in0_1_23: unsigned((21 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((22 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_f0ca8483cb is
  port (
    input_port : in std_logic_vector((21 - 1) downto 0);
    output_port : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_f0ca8483cb;


architecture behavior of reinterpret_f0ca8483cb is
  signal input_port_1_40: signed((21 - 1) downto 0);
  signal output_port_5_5_force: unsigned((21 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_6358c585f1 is
  port (
    a : in std_logic_vector((22 - 1) downto 0);
    b : in std_logic_vector((19 - 1) downto 0);
    s : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_6358c585f1;


architecture behavior of addsub_6358c585f1 is
  signal a_17_32: signed((22 - 1) downto 0);
  signal b_17_35: unsigned((19 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (3 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_91_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_91_20_back: signed((18 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (3 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((23 - 1) downto 0);
  signal cast_69_22: signed((23 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((23 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((18 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(2);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(2);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 2 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 19, 23, 19);
  cast_69_22 <= u2s_cast(b_17_35, 19, 23, 19);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 19, 18, 17);
  op_mem_91_20_front_din <= cast_internal_s_83_3_convert;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_c84451c80b is
  port (
    input_port : in std_logic_vector((22 - 1) downto 0);
    output_port : out std_logic_vector((22 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_c84451c80b;


architecture behavior of reinterpret_c84451c80b is
  signal input_port_1_40: unsigned((22 - 1) downto 0);
  signal output_port_5_5_force: signed((22 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_3013ab8805 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_3013ab8805;


architecture behavior of logical_3013ab8805 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (3 - 1)) of std_logic;
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    '0',
    '0',
    '0');
  signal latency_pipe_5_26_front_din: std_logic;
  signal latency_pipe_5_26_back: std_logic;
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal bit_2_27: std_logic;
  signal fully_2_1_bitnot: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(2);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          latency_pipe_5_26(i) <= latency_pipe_5_26(i-1);
        end loop;
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  bit_2_27 <= d0_1_24 and d1_1_27 and d2_1_30;
  fully_2_1_bitnot <= not bit_2_27;
  latency_pipe_5_26_front_din <= fully_2_1_bitnot;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= std_logic_to_vector(latency_pipe_5_26_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_356a264444 is
  port (
    in0 : in std_logic_vector((21 - 1) downto 0);
    in1 : in std_logic_vector((21 - 1) downto 0);
    in2 : in std_logic_vector((21 - 1) downto 0);
    in3 : in std_logic_vector((21 - 1) downto 0);
    y : out std_logic_vector((84 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_356a264444;


architecture behavior of concat_356a264444 is
  signal in0_1_23: unsigned((21 - 1) downto 0);
  signal in1_1_27: unsigned((21 - 1) downto 0);
  signal in2_1_31: unsigned((21 - 1) downto 0);
  signal in3_1_35: unsigned((21 - 1) downto 0);
  signal y_2_1_concat: unsigned((84 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_43b12feb7d is
  port (
    a : in std_logic_vector((21 - 1) downto 0);
    b : in std_logic_vector((19 - 1) downto 0);
    s : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_43b12feb7d;


architecture behavior of addsub_43b12feb7d is
  signal a_17_32: signed((21 - 1) downto 0);
  signal b_17_35: unsigned((19 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (1 - 1)) of signed((21 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    0 => "000000000000000000000");
  signal op_mem_91_20_front_din: signed((21 - 1) downto 0);
  signal op_mem_91_20_back: signed((21 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (1 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    0 => "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((22 - 1) downto 0);
  signal cast_69_22: signed((22 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((22 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((21 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(0);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(0);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 19, 22, 19);
  cast_69_22 <= u2s_cast(b_17_35, 19, 22, 19);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 19, 21, 18);
  op_mem_91_20_push_front_pop_back_en <= '0';
  cout_mem_92_22_push_front_pop_back_en <= '0';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(cast_internal_s_83_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity scale_97239b8ed2 is
  port (
    ip : in std_logic_vector((20 - 1) downto 0);
    op : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end scale_97239b8ed2;


architecture behavior of scale_97239b8ed2 is
  signal ip_17_23: signed((20 - 1) downto 0);
begin
  ip_17_23 <= std_logic_vector_to_signed(ip);
  op <= signed_to_std_logic_vector(ip_17_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_83820b2faf is
  port (
    in0 : in std_logic_vector((37 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_83820b2faf;


architecture behavior of concat_83820b2faf is
  signal in0_1_23: unsigned((37 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((38 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_db4c53ade5 is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_db4c53ade5;


architecture behavior of reinterpret_db4c53ade5 is
  signal input_port_1_40: signed((37 - 1) downto 0);
  signal output_port_5_5_force: unsigned((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_82254b26db is
  port (
    a : in std_logic_vector((38 - 1) downto 0);
    b : in std_logic_vector((35 - 1) downto 0);
    s : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_82254b26db;


architecture behavior of addsub_82254b26db is
  signal a_17_32: signed((38 - 1) downto 0);
  signal b_17_35: unsigned((35 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (3 - 1)) of signed((19 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "0000000000000000000",
    "0000000000000000000",
    "0000000000000000000");
  signal op_mem_91_20_front_din: signed((19 - 1) downto 0);
  signal op_mem_91_20_back: signed((19 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (3 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((39 - 1) downto 0);
  signal cast_69_22: signed((39 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((39 - 1) downto 0);
  signal cast_internal_s_83_3_convert: signed((19 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(2);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(2);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 2 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 35, 39, 35);
  cast_69_22 <= u2s_cast(b_17_35, 35, 39, 35);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= s2s_cast(internal_s_69_5_addsub, 35, 19, 17);
  op_mem_91_20_front_din <= cast_internal_s_83_3_convert;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_2da6af93c2 is
  port (
    op : out std_logic_vector((35 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_2da6af93c2;


architecture behavior of constant_2da6af93c2 is
begin
  op <= "00000000000000000011111111111111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_620dd01637 is
  port (
    input_port : in std_logic_vector((38 - 1) downto 0);
    output_port : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_620dd01637;


architecture behavior of reinterpret_620dd01637 is
  signal input_port_1_40: unsigned((38 - 1) downto 0);
  signal output_port_5_5_force: signed((38 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_ec14c62a89 is
  port (
    input_port : in std_logic_vector((35 - 1) downto 0);
    output_port : out std_logic_vector((35 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_ec14c62a89;


architecture behavior of reinterpret_ec14c62a89 is
  signal input_port_1_40: unsigned((35 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_5b4829fb41 is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_5b4829fb41;


architecture behavior of reinterpret_5b4829fb41 is
  signal input_port_1_40: unsigned((37 - 1) downto 0);
  signal output_port_5_5_force: signed((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_64530ed2c8 is
  port (
    d : in std_logic_vector((37 - 1) downto 0);
    q : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_64530ed2c8;


architecture behavior of delay_64530ed2c8 is
  signal d_1_22: std_logic_vector((37 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_b28df1ab2e is
  port (
    in0 : in std_logic_vector((36 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_b28df1ab2e;


architecture behavior of concat_b28df1ab2e is
  signal in0_1_23: unsigned((36 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((36 - 1) downto 0);
  signal y_2_1_concat: unsigned((73 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_892b735f0d is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_892b735f0d;


architecture behavior of reinterpret_892b735f0d is
  signal input_port_1_40: unsigned((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_efdf1c3890 is
  port (
    input_port : in std_logic_vector((74 - 1) downto 0);
    output_port : out std_logic_vector((74 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_efdf1c3890;


architecture behavior of reinterpret_efdf1c3890 is
  signal input_port_1_40: unsigned((74 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_56d57d2c92 is
  port (
    in0 : in std_logic_vector((37 - 1) downto 0);
    in1 : in std_logic_vector((37 - 1) downto 0);
    y : out std_logic_vector((74 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_56d57d2c92;


architecture behavior of concat_56d57d2c92 is
  signal in0_1_23: unsigned((37 - 1) downto 0);
  signal in1_1_27: unsigned((37 - 1) downto 0);
  signal y_2_1_concat: unsigned((74 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_4ded11ba54 is
  port (
    a : in std_logic_vector((36 - 1) downto 0);
    b : in std_logic_vector((36 - 1) downto 0);
    s : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_4ded11ba54;


architecture behavior of addsub_4ded11ba54 is
  signal a_17_32: signed((36 - 1) downto 0);
  signal b_17_35: signed((36 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (2 - 1)) of signed((37 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_91_20_front_din: signed((37 - 1) downto 0);
  signal op_mem_91_20_back: signed((37 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (2 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((37 - 1) downto 0);
  signal cast_69_22: signed((37 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((37 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_signed(b);
  op_mem_91_20_back <= op_mem_91_20(1);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(1);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 1 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 34, 37, 34);
  cast_69_22 <= s2s_cast(b_17_35, 34, 37, 34);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  op_mem_91_20_front_din <= internal_s_69_5_addsub;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_8dd4a43ef5 is
  port (
    a : in std_logic_vector((36 - 1) downto 0);
    b : in std_logic_vector((36 - 1) downto 0);
    s : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_8dd4a43ef5;


architecture behavior of addsub_8dd4a43ef5 is
  signal a_17_32: signed((36 - 1) downto 0);
  signal b_17_35: signed((36 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (2 - 1)) of signed((37 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_91_20_front_din: signed((37 - 1) downto 0);
  signal op_mem_91_20_back: signed((37 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (2 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_71_18: signed((37 - 1) downto 0);
  signal cast_71_22: signed((37 - 1) downto 0);
  signal internal_s_71_5_addsub: signed((37 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_signed(b);
  op_mem_91_20_back <= op_mem_91_20(1);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(1);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 1 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_71_18 <= s2s_cast(a_17_32, 34, 37, 34);
  cast_71_22 <= s2s_cast(b_17_35, 34, 37, 34);
  internal_s_71_5_addsub <= cast_71_18 - cast_71_22;
  op_mem_91_20_front_din <= internal_s_71_5_addsub;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mult_f295e5f0f2 is
  port (
    a : in std_logic_vector((18 - 1) downto 0);
    b : in std_logic_vector((18 - 1) downto 0);
    p : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mult_f295e5f0f2;


architecture behavior of mult_f295e5f0f2 is
  signal a_1_22: signed((18 - 1) downto 0);
  signal b_1_25: signed((18 - 1) downto 0);
  type array_type_op_mem_65_20 is array (0 to (2 - 1)) of signed((36 - 1) downto 0);
  signal op_mem_65_20: array_type_op_mem_65_20 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_65_20_front_din: signed((36 - 1) downto 0);
  signal op_mem_65_20_back: signed((36 - 1) downto 0);
  signal op_mem_65_20_push_front_pop_back_en: std_logic;
  signal mult_46_56: signed((36 - 1) downto 0);
begin
  a_1_22 <= std_logic_vector_to_signed(a);
  b_1_25 <= std_logic_vector_to_signed(b);
  op_mem_65_20_back <= op_mem_65_20(1);
  proc_op_mem_65_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_65_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_65_20(i) <= op_mem_65_20(i-1);
        end loop;
        op_mem_65_20(0) <= op_mem_65_20_front_din;
      end if;
    end if;
  end process proc_op_mem_65_20;
  mult_46_56 <= (a_1_22 * b_1_25);
  op_mem_65_20_front_din <= mult_46_56;
  op_mem_65_20_push_front_pop_back_en <= '1';
  p <= signed_to_std_logic_vector(op_mem_65_20_back);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_2d0f74b2c1 is
  port (
    d : in std_logic_vector((37 - 1) downto 0);
    q : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_2d0f74b2c1;


architecture behavior of delay_2d0f74b2c1 is
  signal d_1_22: std_logic_vector((37 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_0cc72cd991 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_0cc72cd991;


architecture behavior of concat_0cc72cd991 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9779a5cf83 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9779a5cf83;


architecture behavior of concat_9779a5cf83 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cda50df78a is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cda50df78a;


architecture behavior of constant_cda50df78a is
begin
  op <= "00";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7eef56098d is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7eef56098d;


architecture behavior of concat_7eef56098d is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_09771002d6 is
  port (
    d : in std_logic_vector((9 - 1) downto 0);
    q : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_09771002d6;


architecture behavior of delay_09771002d6 is
  signal d_1_22: std_logic_vector((9 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000");
  signal op_mem_20_24_front_din: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_pipeline is
    generic (
        old_width   : integer := 16;
        old_bin_pt  : integer := 4;
        old_arith   : integer := xlUnsigned;
        new_width   : integer := 8;
        new_bin_pt  : integer := 2;
        new_arith   : integer := xlUnsigned;
        en_width    : integer := 1;
        en_bin_pt   : integer := 0;
        en_arith    : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow    : integer := xlWrap;
        latency     : integer := 1);
    port (
        din : in std_logic_vector (old_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        result : out std_logic_vector (new_width-1 downto 0));
end convert_pipeline;
architecture behavior of convert_pipeline is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i           : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    constant fp_width : integer := old_width + 2;
    constant fp_bin_pt : integer := old_bin_pt;
    constant fp_arith : integer := old_arith;
    constant q_width : integer := (old_width + 2) + (new_bin_pt - old_bin_pt);
    constant q_bin_pt : integer := new_bin_pt;
    constant q_arith : integer := old_arith;
    signal full_precision_result_in, full_precision_result_out
        : std_logic_vector(fp_width-1 downto 0);
    signal quantized_result_in, quantized_result_out
        : std_logic_vector(q_width-1 downto 0);
    signal result_in : std_logic_vector(new_width-1 downto 0):= (others => '0');
    signal internal_ce : std_logic;
begin
    internal_ce <= ce and en(0);

    fp_result : process (din)
    begin
        full_precision_result_in <= cast(din, old_bin_pt,
                                         fp_width, fp_bin_pt, fp_arith);
    end process;
    latency_fpr : if (latency > 2)
    generate
        reg_fpr : synth_reg
            generic map ( width => fp_width,
                          latency => 1)
            port map (i => full_precision_result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => full_precision_result_out);
    end generate;
    no_latency_fpr : if (latency < 3)
    generate
        full_precision_result_out <= full_precision_result_in;
    end generate;
    xlround_generate : if (quantization = xlRound)
    generate
      xlround_result : process (full_precision_result_out)
      begin
          quantized_result_in <= round_towards_inf(full_precision_result_out,
                                                   fp_width, fp_bin_pt,
                                                   fp_arith, q_width, q_bin_pt,
                                                   q_arith);
      end process;
    end generate;
    xlroundbanker_generate : if (quantization = xlRoundBanker)
    generate
      xlroundbanker_result : process (full_precision_result_out)
      begin
          quantized_result_in <= round_towards_even(full_precision_result_out,
                                                   fp_width, fp_bin_pt,
                                                   fp_arith, q_width, q_bin_pt,
                                                   q_arith);
      end process;
    end generate;
    xltruncate_generate : if (quantization = xlTruncate)
    generate
      xltruncate_result : process (full_precision_result_out)
      begin
          quantized_result_in <= trunc(full_precision_result_out,
                                       fp_width, fp_bin_pt,
                                       fp_arith, q_width, q_bin_pt,
                                       q_arith);
      end process;
    end generate;
    latency_qr : if (latency > 1)
    generate
        reg_qr : synth_reg
            generic map ( width => q_width,
                          latency => 1)
            port map (i => quantized_result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => quantized_result_out);
    end generate;
    no_latency_qr : if (latency < 2)
    generate
        quantized_result_out <= quantized_result_in;
    end generate;
    xlsaturate_generate : if (overflow = xlSaturate)
    generate
      xlsaturate_result : process (quantized_result_out)
      begin
          result_in <= saturation_arith(quantized_result_out, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
      end process;
    end generate;
    xlwrap_generate : if (overflow = xlWrap)
    generate
      xlwrap_result : process (quantized_result_out)
      begin
          result_in <= wrap_arith(quantized_result_out, q_width, q_bin_pt,
                                  q_arith, new_width, new_bin_pt, new_arith);
      end process;
    end generate;
    latency_gt_3 : if (latency > 3)
    generate
        reg_out : synth_reg
            generic map ( width => new_width,
                          latency => latency-2)
            port map (i => result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => result);
    end generate;
    latency_lt_4 : if ((latency < 4) and (latency > 0))
    generate
        reg_out : synth_reg
            generic map ( width => new_width,
                          latency => 1)
            port map (i => result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => result);
    end generate;
    latency0 : if (latency = 0)
    generate
        result <= result_in;
    end generate latency0;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert_pipeline is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din  : in std_logic_vector (din_width-1 downto 0);
        en   : in std_logic_vector (en_width-1 downto 0);
        ce   : in std_logic;
        clr  : in std_logic;
        clk  : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert_pipeline;
architecture behavior of xlconvert_pipeline is
    component convert_pipeline
        generic (
            old_width    : integer := 16;
            old_bin_pt   : integer := 4;
            old_arith    : integer := xlUnsigned;
            new_width    : integer := 8;
            new_bin_pt   : integer := 2;
            new_arith    : integer := xlUnsigned;
            en_width     : integer := 1;
            en_bin_pt    : integer := 0;
            en_arith     : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap;
            latency      : integer := 1);
        port (
            din    : in std_logic_vector (din_width-1 downto 0);
            en     : in std_logic_vector (en_width-1 downto 0);
            ce     : in std_logic;
            clr    : in std_logic;
            clk    : in std_logic;
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
   begin
      convert : convert_pipeline
        generic map (
          old_width   => din_width,
          old_bin_pt  => din_bin_pt,
          old_arith   => din_arith,
          new_width   => dout_width,
          new_bin_pt  => dout_bin_pt,
          new_arith   => dout_arith,
          en_width    => en_width,
          en_bin_pt   => en_bin_pt,
          en_arith    => en_arith,
          quantization => quantization,
          overflow    => overflow,
          latency     => latency)
        port map (
          din => din,
          en => en,
          ce => ce,
          clr => clr,
          clk => clk,
          result => dout);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a7e2bb9e12 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a7e2bb9e12;


architecture behavior of constant_a7e2bb9e12 is
begin
  op <= "01";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4e7d828d94 is
  port (
    d : in std_logic_vector((73 - 1) downto 0);
    q : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4e7d828d94;


architecture behavior of delay_4e7d828d94 is
  signal d_1_22: std_logic_vector((73 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_b6092ad150 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_b6092ad150;


architecture behavior of delay_b6092ad150 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_206b7f76d8 is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_206b7f76d8;


architecture behavior of negate_206b7f76d8 is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (1 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    0 => "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(0);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  internal_ip_40_3_convert <= std_logic_vector_to_signed(convert_type(signed_to_std_logic_vector(internal_ip_join_30_1), 19, 17, xlSigned, 18, 17, xlSigned, xlTruncate, xlSaturate));
  op_mem_48_20_front_din <= internal_ip_40_3_convert;
  op_mem_48_20_push_front_pop_back_en <= '1';
  op <= signed_to_std_logic_vector(op_mem_48_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_bc64561e19 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_bc64561e19;


architecture behavior of mux_bc64561e19 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_7097453b2c is
  port (
    d : in std_logic_vector((73 - 1) downto 0);
    q : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_7097453b2c;


architecture behavior of delay_7097453b2c is
  signal d_1_22: std_logic_vector((73 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlpassthrough is
    generic (
        din_width    : integer := 16;
        dout_width   : integer := 16
        );
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlpassthrough;
architecture passthrough_arch of xlpassthrough is
begin
  dout <= din;
end passthrough_arch;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xldpram_fft_core is
  generic (
    core_name0: string := "";
    c_width_a: integer := 13;
    c_address_width_a: integer := 4;
    c_width_b: integer := 13;
    c_address_width_b: integer := 4;
    c_has_sinita: integer := 0;
    c_has_sinitb: integer := 0;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width_a - 1 downto 0);
    addra: in std_logic_vector(c_address_width_a - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    a_ce: in std_logic;
    a_clk: in std_logic;
    rsta: in std_logic_vector(0 downto 0) := (others => '0');
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    douta: out std_logic_vector(c_width_a - 1 downto 0);
    dinb: in std_logic_vector(c_width_b - 1 downto 0);
    addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
    web: in std_logic_vector(0 downto 0);
    b_ce: in std_logic;
    b_clk: in std_logic;
    rstb: in std_logic_vector(0 downto 0) := (others => '0');
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    doutb: out std_logic_vector(c_width_b - 1 downto 0)
  );
end xldpram_fft_core;
architecture behavior of xldpram_fft_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;

  signal core_addra: std_logic_vector(c_address_width_a - 1 downto 0);
  signal core_addrb: std_logic_vector(c_address_width_b - 1 downto 0);
  signal core_dina, core_douta, dly_douta:
    std_logic_vector(c_width_a - 1 downto 0);
  signal core_dinb, core_doutb, dly_doutb:
    std_logic_vector(c_width_b - 1 downto 0);
  signal core_wea, core_web: std_logic;
  signal core_a_ce, core_b_ce: std_logic;
  signal sinita, sinitb: std_logic;

  component bmg_72_c1a8b20e2e422729
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_c1a8b20e2e422729:
    component is true;
  attribute fpga_dont_touch of bmg_72_c1a8b20e2e422729:
    component is "true";
  attribute box_type of bmg_72_c1a8b20e2e422729:
    component  is "black_box";
  component bmg_72_9f585cf1e3329833
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_9f585cf1e3329833:
    component is true;
  attribute fpga_dont_touch of bmg_72_9f585cf1e3329833:
    component is "true";
  attribute box_type of bmg_72_9f585cf1e3329833:
    component  is "black_box";
  component bmg_72_488bc588e4c66edf
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_488bc588e4c66edf:
    component is true;
  attribute fpga_dont_touch of bmg_72_488bc588e4c66edf:
    component is "true";
  attribute box_type of bmg_72_488bc588e4c66edf:
    component  is "black_box";
  component bmg_72_53d3a85261e207bb
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_53d3a85261e207bb:
    component is true;
  attribute fpga_dont_touch of bmg_72_53d3a85261e207bb:
    component is "true";
  attribute box_type of bmg_72_53d3a85261e207bb:
    component  is "black_box";
begin
  core_addra <= addra;
  core_dina <= dina;
  douta <= dly_douta;
  core_wea <= wea(0);
  core_a_ce <= a_ce and ena(0);
  sinita <= rsta(0) and a_ce;

  core_addrb <= addrb;
  core_dinb <= dinb;
  doutb <= dly_doutb;
  core_web <= web(0);
  core_b_ce <= b_ce and enb(0);
  sinitb <= rstb(0) and b_ce;
  comp0: if ((core_name0 = "bmg_72_c1a8b20e2e422729")) generate
    core_instance0: bmg_72_c1a8b20e2e422729
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_9f585cf1e3329833")) generate
    core_instance1: bmg_72_9f585cf1e3329833
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp2: if ((core_name0 = "bmg_72_488bc588e4c66edf")) generate
    core_instance2: bmg_72_488bc588e4c66edf
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp3: if ((core_name0 = "bmg_72_53d3a85261e207bb")) generate
    core_instance3: bmg_72_53d3a85261e207bb
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  latency_test: if (latency > 2) generate
    regA: synth_reg
      generic map (
        width => c_width_a,
        latency => latency - 2
      )
      port map (
        i => core_douta,
        ce => core_a_ce,
        clr => '0',
        clk => a_clk,
        o => dly_douta
      );
    regB: synth_reg
      generic map (
        width => c_width_b,
        latency => latency - 2
      )
      port map (
        i => core_doutb,
        ce => core_b_ce,
        clr => '0',
        clk => b_clk,
        o => dly_doutb
      );
  end generate;
  latency1: if (latency <= 2) generate
    dly_douta <= core_douta;
    dly_doutb <= core_doutb;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_95b0f967bc is
  port (
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_95b0f967bc;


architecture behavior of constant_95b0f967bc is
begin
  op <= "000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_cfdc93535e is
  port (
    in0 : in std_logic_vector((40 - 1) downto 0);
    in1 : in std_logic_vector((40 - 1) downto 0);
    y : out std_logic_vector((80 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_cfdc93535e;


architecture behavior of concat_cfdc93535e is
  signal in0_1_23: unsigned((40 - 1) downto 0);
  signal in1_1_27: unsigned((40 - 1) downto 0);
  signal y_2_1_concat: unsigned((80 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_86d5838e9c is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((84 - 1) downto 0);
    d1 : in std_logic_vector((84 - 1) downto 0);
    y : out std_logic_vector((84 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_86d5838e9c;


architecture behavior of mux_86d5838e9c is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((84 - 1) downto 0);
  signal d1_1_27: std_logic_vector((84 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((84 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    "000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((84 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((84 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((84 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_faa52967c8 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_faa52967c8;


architecture behavior of delay_faa52967c8 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (8 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(7);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 7 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_67ad97ca70 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_67ad97ca70;


architecture behavior of constant_67ad97ca70 is
begin
  op <= "0001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_145086465d is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_145086465d;


architecture behavior of constant_145086465d is
begin
  op <= "1000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_4d3cfceaf4 is
  port (
    a : in std_logic_vector((4 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_4d3cfceaf4;


architecture behavior of relational_4d3cfceaf4 is
  signal a_1_31: unsigned((4 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e774b32dc9 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e774b32dc9;


architecture behavior of concat_e774b32dc9 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_811dd91a3d is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((10 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_811dd91a3d;


architecture behavior of concat_811dd91a3d is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((10 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4fd36a24a3 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4fd36a24a3;


architecture behavior of concat_4fd36a24a3 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_cf4f99539f is
  port (
    d : in std_logic_vector((10 - 1) downto 0);
    q : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_cf4f99539f;


architecture behavior of delay_cf4f99539f is
  signal d_1_22: std_logic_vector((10 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000000000");
  signal op_mem_20_24_front_din: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a1c496ea88 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a1c496ea88;


architecture behavior of constant_a1c496ea88 is
begin
  op <= "001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_822933f89b is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_822933f89b;


architecture behavior of constant_822933f89b is
begin
  op <= "000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_469094441c is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_469094441c;


architecture behavior of constant_469094441c is
begin
  op <= "100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_8fc7f5539b is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_8fc7f5539b;


architecture behavior of relational_8fc7f5539b is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_47b317dab6 is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_47b317dab6;


architecture behavior of relational_47b317dab6 is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0fa71d0d3 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    in10 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0fa71d0d3;


architecture behavior of concat_a0fa71d0d3 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal in10_1_63: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  in10_1_63 <= std_logic_vector_to_unsigned(in10);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59) & unsigned_to_std_logic_vector(in10_1_63));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9769d05421 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((11 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9769d05421;


architecture behavior of concat_9769d05421 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((11 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7ad1e33701 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((10 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7ad1e33701;


architecture behavior of concat_7ad1e33701 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((10 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_49cb1051e0 is
  port (
    d : in std_logic_vector((11 - 1) downto 0);
    q : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_49cb1051e0;


architecture behavior of delay_49cb1051e0 is
  signal d_1_22: std_logic_vector((11 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000000000");
  signal op_mem_20_24_front_din: std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_38898c80c0 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_38898c80c0;


architecture behavior of delay_38898c80c0 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8ddc079e9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8ddc079e9;


architecture behavior of constant_e8ddc079e9 is
begin
  op <= "10";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5f1eb17108 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5f1eb17108;


architecture behavior of relational_5f1eb17108 is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_f9928864ea is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_f9928864ea;


architecture behavior of relational_f9928864ea is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ef66525e56 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    in10 : in std_logic_vector((1 - 1) downto 0);
    in11 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ef66525e56;


architecture behavior of concat_ef66525e56 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal in10_1_63: unsigned((1 - 1) downto 0);
  signal in11_1_68: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  in10_1_63 <= std_logic_vector_to_unsigned(in10);
  in11_1_68 <= std_logic_vector_to_unsigned(in11);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59) & unsigned_to_std_logic_vector(in10_1_63) & unsigned_to_std_logic_vector(in11_1_68));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_118109a960 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_118109a960;


architecture behavior of concat_118109a960 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((12 - 1) downto 0);
  signal y_2_1_concat: unsigned((13 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_8503582fb5 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((11 - 1) downto 0);
    y : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_8503582fb5;


architecture behavior of concat_8503582fb5 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((11 - 1) downto 0);
  signal y_2_1_concat: unsigned((13 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_87cc993d41 is
  port (
    d : in std_logic_vector((12 - 1) downto 0);
    q : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_87cc993d41;


architecture behavior of delay_87cc993d41 is
  signal d_1_22: std_logic_vector((12 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_9b03e3d644 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_9b03e3d644;


architecture behavior of counter_9b03e3d644 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((1 - 1) downto 0) := "0";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((2 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("1");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_894f23b88c is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_894f23b88c;


architecture behavior of negate_894f23b88c is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (4 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(3);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop 
          op_mem_48_20(i) <= op_mem_48_20(i-1);
        end loop;
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  internal_ip_40_3_convert <= std_logic_vector_to_signed(convert_type(signed_to_std_logic_vector(internal_ip_join_30_1), 19, 17, xlSigned, 18, 17, xlSigned, xlTruncate, xlSaturate));
  op_mem_48_20_front_din <= internal_ip_40_3_convert;
  op_mem_48_20_push_front_pop_back_en <= '1';
  op <= signed_to_std_logic_vector(op_mem_48_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_8f386731a6 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_8f386731a6;


architecture behavior of counter_8f386731a6 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((12 - 1) downto 0) := "000000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((13 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4c85700954 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4c85700954;


architecture behavior of delay_4c85700954 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (10 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(9);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 9 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_5b3ce5f2ae is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_5b3ce5f2ae;


architecture behavior of delay_5b3ce5f2ae is
  signal d_1_22: std_logic_vector((1 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (6 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0",
    "0",
    "0",
    "0",
    "0",
    "0");
  signal op_mem_20_24_front_din: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(5);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4217913c13 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4217913c13;


architecture behavior of delay_4217913c13 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (6 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(5);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_c462a80bee is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_c462a80bee;


architecture behavior of delay_c462a80bee is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_328e8ebbb5 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_328e8ebbb5;


architecture behavior of delay_328e8ebbb5 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_30e9ca90db is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_30e9ca90db;


architecture behavior of mux_30e9ca90db is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (7 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(6);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 6 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_181e58d842 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_181e58d842;


architecture behavior of mux_181e58d842 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7c91b1b314 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7c91b1b314;


architecture behavior of constant_7c91b1b314 is
begin
  op <= "000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd28b32bf8 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd28b32bf8;


architecture behavior of constant_fd28b32bf8 is
begin
  op <= "000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e054d850c5 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e054d850c5;


architecture behavior of constant_e054d850c5 is
begin
  op <= "100000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_d36fe12c1c is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_d36fe12c1c;


architecture behavior of relational_d36fe12c1c is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_acb3c05dd0 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_acb3c05dd0;


architecture behavior of relational_acb3c05dd0 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e6f5ee726b is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e6f5ee726b;


architecture behavior of concat_e6f5ee726b is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((2 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4a9a9a25a3 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4a9a9a25a3;


architecture behavior of concat_4a9a9a25a3 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((2 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_6160d7387c is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_6160d7387c;


architecture behavior of concat_6160d7387c is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4ce33ca7e7 is
  port (
    d : in std_logic_vector((2 - 1) downto 0);
    q : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4ce33ca7e7;


architecture behavior of delay_4ce33ca7e7 is
  signal d_1_22: std_logic_vector((2 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00");
  signal op_mem_20_24_front_din: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldpram_dist_fft_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    addr_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width - 1 downto 0);
    addra: in std_logic_vector(addr_width - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    a_ce: in std_logic;
    a_clk: in std_logic;
    douta: out std_logic_vector(c_width - 1 downto 0);
    addrb: in std_logic_vector(addr_width - 1 downto 0);
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    b_ce: in std_logic;
    b_clk: in std_logic;
    doutb: out std_logic_vector(c_width - 1 downto 0)
  );
end xldpram_dist_fft_core ;
architecture behavior of xldpram_dist_fft_core is
  component synth_reg is
    generic (
      width: integer := 8;
      latency: integer := 1
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  constant num_extra_addr_bits: integer := (c_address_width - addr_width);
  signal core_addra, core_addrb: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_in, core_douta, core_doutb: std_logic_vector(c_width - 1 downto 0);
  signal reg_douta, reg_doutb: std_logic_vector(c_width - 1 downto 0);
  signal core_we: std_logic_vector(0 downto 0);
  signal core_cea, core_ceb: std_logic;
  component dmg_72_505931c5b3ea228e
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_505931c5b3ea228e:
    component is true;
  attribute fpga_dont_touch of dmg_72_505931c5b3ea228e:
    component is "true";
  attribute box_type of dmg_72_505931c5b3ea228e:
    component  is "black_box";
  component dmg_72_d20b02a9f8239c7a
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_d20b02a9f8239c7a:
    component is true;
  attribute fpga_dont_touch of dmg_72_d20b02a9f8239c7a:
    component is "true";
  attribute box_type of dmg_72_d20b02a9f8239c7a:
    component  is "black_box";
  component dmg_72_efdf1b1b05926829
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_efdf1b1b05926829:
    component is true;
  attribute fpga_dont_touch of dmg_72_efdf1b1b05926829:
    component is "true";
  attribute box_type of dmg_72_efdf1b1b05926829:
    component  is "black_box";
  component dmg_72_1c323e86177437db
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_1c323e86177437db:
    component is true;
  attribute fpga_dont_touch of dmg_72_1c323e86177437db:
    component is "true";
  attribute box_type of dmg_72_1c323e86177437db:
    component  is "black_box";
begin
  need_to_pad_addr : if num_extra_addr_bits > 0 generate
      core_addra(c_address_width - 1 downto addr_width) <= (others => '0');
      core_addra(addr_width - 1 downto 0) <= addra;
      core_addrb(c_address_width - 1 downto addr_width) <= (others => '0');
      core_addrb(addr_width - 1 downto 0) <= addrb;
  end generate;
  no_need_to_pad_addr: if num_extra_addr_bits = 0 generate
    core_addra <= addra;
    core_addrb <= addrb;
  end generate;
  douta <= reg_douta;
  doutb <= reg_doutb;
  core_cea <= a_ce and ena(0);
  core_ceb <= b_ce and enb(0);
  core_we(0) <= wea(0) and core_cea;
  registered_dpram : if latency > 0 generate
    output_rega: synth_reg
      generic map (
        width   => c_width,
        latency => latency
      )
      port map (
        i   => core_douta,
        ce  => core_cea,
        clr => '0',
        clk => a_clk,
        o   => reg_douta
      );
    output_regb: synth_reg
      generic map (
        width   => c_width,
        latency => latency
      )
      port map (
        i   => core_doutb,
        ce  => core_ceb,
        clr => '0',
        clk => b_clk,
        o   => reg_doutb
      );
  end generate;
  nonregistered_ram : if latency = 0 generate
    reg_douta <= core_douta;
    reg_doutb <= core_doutb;
  end generate;
  comp0: if ((core_name0 = "dmg_72_505931c5b3ea228e")) generate
    core_instance0: dmg_72_505931c5b3ea228e
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "dmg_72_d20b02a9f8239c7a")) generate
    core_instance1: dmg_72_d20b02a9f8239c7a
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp2: if ((core_name0 = "dmg_72_efdf1b1b05926829")) generate
    core_instance2: dmg_72_efdf1b1b05926829
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp3: if ((core_name0 = "dmg_72_1c323e86177437db")) generate
    core_instance3: dmg_72_1c323e86177437db
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_118598964d is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_118598964d;


architecture behavior of constant_118598964d is
begin
  op <= "00000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a3923dd146 is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a3923dd146;


architecture behavior of constant_a3923dd146 is
begin
  op <= "00000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0604807f72 is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0604807f72;


architecture behavior of constant_0604807f72 is
begin
  op <= "10000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2147430058 is
  port (
    a : in std_logic_vector((11 - 1) downto 0);
    b : in std_logic_vector((11 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2147430058;


architecture behavior of relational_2147430058 is
  signal a_1_31: unsigned((11 - 1) downto 0);
  signal b_1_34: unsigned((11 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_b4b277ae0f is
  port (
    a : in std_logic_vector((11 - 1) downto 0);
    b : in std_logic_vector((11 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_b4b277ae0f;


architecture behavior of relational_b4b277ae0f is
  signal a_1_31: unsigned((11 - 1) downto 0);
  signal b_1_34: unsigned((11 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_452c4d3410 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_452c4d3410;


architecture behavior of concat_452c4d3410 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_949f038a6d is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_949f038a6d;


architecture behavior of concat_949f038a6d is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_54d5af2115 is
  port (
    d : in std_logic_vector((3 - 1) downto 0);
    q : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_54d5af2115;


architecture behavior of delay_54d5af2115 is
  signal d_1_22: std_logic_vector((3 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000");
  signal op_mem_20_24_front_din: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_f1ac4bddff is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_f1ac4bddff;


architecture behavior of constant_f1ac4bddff is
begin
  op <= "0000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_498bc68c14 is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_498bc68c14;


architecture behavior of constant_498bc68c14 is
begin
  op <= "0000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fbc2f0cce1 is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fbc2f0cce1;


architecture behavior of constant_fbc2f0cce1 is
begin
  op <= "1000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_0ffd72e037 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_0ffd72e037;


architecture behavior of relational_0ffd72e037 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_f6702ea2f7 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_f6702ea2f7;


architecture behavior of relational_f6702ea2f7 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_cf540617d5 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_cf540617d5;


architecture behavior of concat_cf540617d5 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_8f12c32de0 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_8f12c32de0;


architecture behavior of concat_8f12c32de0 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4ca77626c8 is
  port (
    d : in std_logic_vector((4 - 1) downto 0);
    q : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4ca77626c8;


architecture behavior of delay_4ca77626c8 is
  signal d_1_22: std_logic_vector((4 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000");
  signal op_mem_20_24_front_din: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b4ec9de7d1 is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b4ec9de7d1;


architecture behavior of constant_b4ec9de7d1 is
begin
  op <= "000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd85eb7067 is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd85eb7067;


architecture behavior of constant_fd85eb7067 is
begin
  op <= "000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4a391b9a0e is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4a391b9a0e;


architecture behavior of constant_4a391b9a0e is
begin
  op <= "100000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6c3ee657fa is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6c3ee657fa;


architecture behavior of relational_6c3ee657fa is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_78eac2928d is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_78eac2928d;


architecture behavior of relational_78eac2928d is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2b3acb49f4 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2b3acb49f4;


architecture behavior of concat_2b3acb49f4 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ac785d9b37 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ac785d9b37;


architecture behavior of concat_ac785d9b37 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ae3f02567e is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ae3f02567e;


architecture behavior of concat_ae3f02567e is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_b096bcf164 is
  port (
    d : in std_logic_vector((5 - 1) downto 0);
    q : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_b096bcf164;


architecture behavior of delay_b096bcf164 is
  signal d_1_22: std_logic_vector((5 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000");
  signal op_mem_20_24_front_din: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b437b02512 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b437b02512;


architecture behavior of constant_b437b02512 is
begin
  op <= "00000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_91ef1678ca is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_91ef1678ca;


architecture behavior of constant_91ef1678ca is
begin
  op <= "00000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8aae5d3bb is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8aae5d3bb;


architecture behavior of constant_e8aae5d3bb is
begin
  op <= "10000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_54048c8b02 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54048c8b02;


architecture behavior of relational_54048c8b02 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_16235eb2bf is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_16235eb2bf;


architecture behavior of relational_16235eb2bf is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2dc093ca7a is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2dc093ca7a;


architecture behavior of concat_2dc093ca7a is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c6a9b6687e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c6a9b6687e;


architecture behavior of concat_c6a9b6687e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_75261c7c53 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_75261c7c53;


architecture behavior of concat_75261c7c53 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0b18d34058 is
  port (
    d : in std_logic_vector((6 - 1) downto 0);
    q : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0b18d34058;


architecture behavior of delay_0b18d34058 is
  signal d_1_22: std_logic_vector((6 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000");
  signal op_mem_20_24_front_din: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_fft_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_fft_core ;
architecture behavior of xlsprom_fft_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_ce, sinit: std_logic;
  component bmg_72_eb304381eda4ae1e
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_eb304381eda4ae1e:
    component is true;
  attribute fpga_dont_touch of bmg_72_eb304381eda4ae1e:
    component is "true";
  attribute box_type of bmg_72_eb304381eda4ae1e:
    component  is "black_box";
  component bmg_72_6711bf92f3a48934
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_6711bf92f3a48934:
    component is true;
  attribute fpga_dont_touch of bmg_72_6711bf92f3a48934:
    component is "true";
  attribute box_type of bmg_72_6711bf92f3a48934:
    component  is "black_box";
  component bmg_72_070de696ab472038
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_070de696ab472038:
    component is true;
  attribute fpga_dont_touch of bmg_72_070de696ab472038:
    component is "true";
  attribute box_type of bmg_72_070de696ab472038:
    component  is "black_box";
begin
  core_addr <= addr;
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_eb304381eda4ae1e")) generate
    core_instance0: bmg_72_eb304381eda4ae1e
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp1: if ((core_name0 = "bmg_72_6711bf92f3a48934")) generate
    core_instance1: bmg_72_6711bf92f3a48934
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp2: if ((core_name0 = "bmg_72_070de696ab472038")) generate
    core_instance2: bmg_72_070de696ab472038
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_1: if (latency <= 1) generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_180df391de is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_180df391de;


architecture behavior of constant_180df391de is
begin
  op <= "0000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7244cd602b is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7244cd602b;


architecture behavior of constant_7244cd602b is
begin
  op <= "0000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7b07120b87 is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7b07120b87;


architecture behavior of constant_7b07120b87 is
begin
  op <= "1000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9a3978c602 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9a3978c602;


architecture behavior of relational_9a3978c602 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_23065a6aa3 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_23065a6aa3;


architecture behavior of relational_23065a6aa3 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_eb5f1ca7f9 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_eb5f1ca7f9;


architecture behavior of concat_eb5f1ca7f9 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_83e473517e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_83e473517e;


architecture behavior of concat_83e473517e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((7 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_dc245eb1d2 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_dc245eb1d2;


architecture behavior of concat_dc245eb1d2 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_9066adfc41 is
  port (
    d : in std_logic_vector((7 - 1) downto 0);
    q : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_9066adfc41;


architecture behavior of delay_9066adfc41 is
  signal d_1_22: std_logic_vector((7 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000000");
  signal op_mem_20_24_front_din: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a267c870be is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a267c870be;


architecture behavior of constant_a267c870be is
begin
  op <= "000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7ea0f2fff7 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7ea0f2fff7;


architecture behavior of constant_7ea0f2fff7 is
begin
  op <= "000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_961b61f8a1 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_961b61f8a1;


architecture behavior of constant_961b61f8a1 is
begin
  op <= "100000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_931d61fb72 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_931d61fb72;


architecture behavior of relational_931d61fb72 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_fe487ce1c7 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_fe487ce1c7;


architecture behavior of relational_fe487ce1c7 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7673b9b993 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7673b9b993;


architecture behavior of concat_7673b9b993 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_1ece14600f is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_1ece14600f;


architecture behavior of concat_1ece14600f is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_f62149b02a is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_f62149b02a;


architecture behavior of concat_f62149b02a is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((7 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_ebec135d8a is
  port (
    d : in std_logic_vector((8 - 1) downto 0);
    q : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_ebec135d8a;


architecture behavior of delay_ebec135d8a is
  signal d_1_22: std_logic_vector((8 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000000");
  signal op_mem_20_24_front_din: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_3a3620b5a6 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_3a3620b5a6;


architecture behavior of delay_3a3620b5a6 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (16 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(15);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 15 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_582a3706dd is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_582a3706dd;


architecture behavior of constant_582a3706dd is
begin
  op <= "00001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fe72737ca0 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fe72737ca0;


architecture behavior of constant_fe72737ca0 is
begin
  op <= "00000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_ef0e2e5fc6 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_ef0e2e5fc6;


architecture behavior of constant_ef0e2e5fc6 is
begin
  op <= "10000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9ece3c8c4e is
  port (
    a : in std_logic_vector((5 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9ece3c8c4e;


architecture behavior of relational_9ece3c8c4e is
  signal a_1_31: unsigned((5 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_dc5bc996c9 is
  port (
    a : in std_logic_vector((5 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_dc5bc996c9;


architecture behavior of relational_dc5bc996c9 is
  signal a_1_31: unsigned((5 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/delay0"

entity delay0_entity_4675455b89 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_4675455b89;

architecture structural of delay0_entity_4675455b89 is
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  reinterpret_out_output_port_net_x0 <= din;
  dout <= ram_data_out_net_x0;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 4092,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_ed810b6704650710",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_77dc1780892a0930",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      data_in => reinterpret_out_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/add_even_real/a_debus"

entity a_debus_entity_459b56afaf is
  port (
    bus_in: in std_logic_vector(17 downto 0); 
    msb_lsb_out1: out std_logic_vector(17 downto 0)
  );
end a_debus_entity_459b56afaf;

architecture structural of a_debus_entity_459b56afaf is
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x0 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 18,
      y_width => 18
    )
    port map (
      x => reinterpret2_output_port_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/add_even_real/op_bussify"

entity op_bussify_entity_a0c10d7209 is
  port (
    in1: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(18 downto 0)
  );
end op_bussify_entity_a0c10d7209;

architecture structural of op_bussify_entity_a0c10d7209 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/add_even_real"

entity add_even_real_entity_d02be0cdd9 is
  port (
    a: in std_logic_vector(17 downto 0); 
    b: in std_logic_vector(17 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(18 downto 0)
  );
end add_even_real_entity_d02be0cdd9;

architecture structural of add_even_real_entity_d02be0cdd9 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x2: std_logic;
  signal clk_1_sg_x2: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x2 <= a;
  reinterpret2_output_port_net_x3 <= b;
  ce_1_sg_x2 <= ce_1;
  clk_1_sg_x2 <= clk_1;
  dout <= reinterpret1_output_port_net_x3;

  a_debus_459b56afaf: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret2_output_port_net_x2,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_59920783799a8e86",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x2,
      clk => clk_1_sg_x2,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  b_debus_571db2539a: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret2_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  op_bussify_a0c10d7209: entity work.op_bussify_entity_a0c10d7209
    port map (
      in1 => addsub1_s_net_x0,
      bus_out => reinterpret1_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_convert/bussify"

entity bussify_entity_1d06622102 is
  port (
    in1: in std_logic_vector(17 downto 0); 
    in2: in std_logic_vector(17 downto 0); 
    in3: in std_logic_vector(17 downto 0); 
    in4: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(71 downto 0)
  );
end bussify_entity_1d06622102;

architecture structural of bussify_entity_1d06622102 is
  signal adder_s_net_x3: std_logic_vector(17 downto 0);
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(17 downto 0);

begin
  adder_s_net_x3 <= in1;
  adder_s_net_x4 <= in2;
  adder_s_net_x5 <= in3;
  adder_s_net_x6 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_a246e373e7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x3,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x4,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x5,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x6,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_convert/conv1"

entity conv1_entity_9b4d843cb7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(18 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end conv1_entity_9b4d843cb7;

architecture structural of conv1_entity_9b4d843cb7 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x4: std_logic;
  signal clk_1_sg_x4: std_logic;
  signal concat_y_net: std_logic_vector(19 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(19 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(18 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x4 <= ce_1;
  clk_1_sg_x4 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.addsub_f4186754a0
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 19,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_504cae28bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_convert/debus"

entity debus_entity_3f078924c3 is
  port (
    bus_in: in std_logic_vector(75 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out4: out std_logic_vector(18 downto 0); 
    out2: out std_logic_vector(18 downto 0); 
    out3: out std_logic_vector(18 downto 0)
  );
end debus_entity_3f078924c3;

architecture structural of debus_entity_3f078924c3 is
  signal concatenate_y_net_x0: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);
  signal slice3_y_net: std_logic_vector(18 downto 0);
  signal slice4_y_net: std_logic_vector(18 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x1;
  msb_out4 <= reinterpret4_output_port_net_x1;
  out2 <= reinterpret2_output_port_net_x1;
  out3 <= reinterpret3_output_port_net_x1;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x1
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x1
    );

  reinterpret3: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x1
    );

  reinterpret4: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 38,
      new_msb => 56,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 57,
      new_msb => 75,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_convert"

entity bus_convert_entity_6fcb7792a1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(71 downto 0)
  );
end bus_convert_entity_6fcb7792a1;

architecture structural of bus_convert_entity_6fcb7792a1 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal ce_1_sg_x8: std_logic;
  signal clk_1_sg_x8: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x8 <= ce_1;
  clk_1_sg_x8 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_1d06622102: entity work.bussify_entity_1d06622102
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_9b4d843cb7: entity work.conv1_entity_9b4d843cb7
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_77aca7cbad: entity work.conv1_entity_9b4d843cb7
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_4f821fbbd8: entity work.conv1_entity_9b4d843cb7
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_44c25e363b: entity work.conv1_entity_9b4d843cb7
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_3f078924c3: entity work.debus_entity_3f078924c3
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_expand"

entity bus_expand_entity_26ad604baf is
  port (
    bus_in: in std_logic_vector(71 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out4: out std_logic_vector(17 downto 0); 
    out2: out std_logic_vector(17 downto 0); 
    out3: out std_logic_vector(17 downto 0)
  );
end bus_expand_entity_26ad604baf;

architecture structural of bus_expand_entity_26ad604baf is
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);
  signal slice3_y_net: std_logic_vector(17 downto 0);
  signal slice4_y_net: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x4 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 53,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 54,
      new_msb => 71,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_expand_a"

entity bus_expand_a_entity_e0cf78c6cc is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out2: out std_logic_vector(17 downto 0)
  );
end bus_expand_a_entity_e0cf78c6cc;

architecture structural of bus_expand_a_entity_e0cf78c6cc is
  signal reinterpret1_output_port_net_x6: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);

begin
  reinterpret_out_output_port_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x6;
  msb_out2 <= reinterpret2_output_port_net_x3;

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x6
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x3
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret_out_output_port_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret_out_output_port_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_scale/bussify"

entity bussify_entity_5c7818bd70 is
  port (
    in1: in std_logic_vector(18 downto 0); 
    in2: in std_logic_vector(18 downto 0); 
    in3: in std_logic_vector(18 downto 0); 
    in4: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(75 downto 0)
  );
end bussify_entity_5c7818bd70;

architecture structural of bussify_entity_5c7818bd70 is
  signal concatenate_y_net_x3: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(18 downto 0);
  signal scale1_op_net_x0: std_logic_vector(18 downto 0);
  signal scale2_op_net_x0: std_logic_vector(18 downto 0);
  signal scale3_op_net_x0: std_logic_vector(18 downto 0);
  signal scale4_op_net_x0: std_logic_vector(18 downto 0);

begin
  scale1_op_net_x0 <= in1;
  scale2_op_net_x0 <= in2;
  scale3_op_net_x0 <= in3;
  scale4_op_net_x0 <= in4;
  bus_out <= concatenate_y_net_x3;

  concatenate: entity work.concat_2aea51ccde
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x3
    );

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale1_op_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale2_op_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale3_op_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale4_op_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_scale/debus"

entity debus_entity_8ef01a3c6c is
  port (
    bus_in: in std_logic_vector(75 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out4: out std_logic_vector(18 downto 0); 
    out2: out std_logic_vector(18 downto 0); 
    out3: out std_logic_vector(18 downto 0)
  );
end debus_entity_8ef01a3c6c;

architecture structural of debus_entity_8ef01a3c6c is
  signal concat_y_net_x0: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);
  signal slice3_y_net: std_logic_vector(18 downto 0);
  signal slice4_y_net: std_logic_vector(18 downto 0);

begin
  concat_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 38,
      new_msb => 56,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 57,
      new_msb => 75,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/bus_scale"

entity bus_scale_entity_472dd14792 is
  port (
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(75 downto 0)
  );
end bus_scale_entity_472dd14792;

architecture structural of bus_scale_entity_472dd14792 is
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal scale1_op_net_x0: std_logic_vector(18 downto 0);
  signal scale2_op_net_x0: std_logic_vector(18 downto 0);
  signal scale3_op_net_x0: std_logic_vector(18 downto 0);
  signal scale4_op_net_x0: std_logic_vector(18 downto 0);

begin
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x4;

  bussify_5c7818bd70: entity work.bussify_entity_5c7818bd70
    port map (
      in1 => scale1_op_net_x0,
      in2 => scale2_op_net_x0,
      in3 => scale3_op_net_x0,
      in4 => scale4_op_net_x0,
      bus_out => concatenate_y_net_x4
    );

  debus_8ef01a3c6c: entity work.debus_entity_8ef01a3c6c
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  scale1: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret4_output_port_net_x0,
      op => scale1_op_net_x0
    );

  scale2: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret3_output_port_net_x0,
      op => scale2_op_net_x0
    );

  scale3: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret2_output_port_net_x0,
      op => scale3_op_net_x0
    );

  scale4: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret1_output_port_net_x0,
      op => scale4_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/munge_a/join"

entity join_entity_dce4ac7e98 is
  port (
    in1: in std_logic_vector(17 downto 0); 
    in2: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end join_entity_dce4ac7e98;

architecture structural of join_entity_dce4ac7e98 is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x1 <= in1;
  reinterpret1_output_port_net_x1 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret1_output_port_net_x1,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/munge_a"

entity munge_a_entity_40c03aaddb is
  port (
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end munge_a_entity_40c03aaddb;

architecture structural of munge_a_entity_40c03aaddb is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal mux0_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(35 downto 0);

begin
  mux0_y_net_x0 <= din;
  dout <= reinterpret_out_output_port_net_x1;

  join_dce4ac7e98: entity work.join_entity_dce4ac7e98
    port map (
      in1 => reinterpret2_output_port_net_x2,
      in2 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x0
    );

  reinterpret: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux0_y_net_x0,
      output_port => reinterpret_output_port_net_x0
    );

  reinterpret_out: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x0,
      output_port => reinterpret_out_output_port_net_x1
    );

  split_5783538a3a: entity work.bus_expand_a_entity_e0cf78c6cc
    port map (
      bus_in => reinterpret_output_port_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/ri_to_c"

entity ri_to_c_entity_2b066e56b4 is
  port (
    im: in std_logic_vector(17 downto 0); 
    re: in std_logic_vector(17 downto 0); 
    c: out std_logic_vector(35 downto 0)
  );
end ri_to_c_entity_2b066e56b4;

architecture structural of ri_to_c_entity_2b066e56b4 is
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal force_im_output_port_net: std_logic_vector(17 downto 0);
  signal force_re_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x1 <= im;
  reinterpret4_output_port_net_x1 <= re;
  c <= concat_y_net_x1;

  concat: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x1
    );

  force_im: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x1,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0/sub_even_imag"

entity sub_even_imag_entity_77ffaad0ab is
  port (
    a: in std_logic_vector(17 downto 0); 
    b: in std_logic_vector(17 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(18 downto 0)
  );
end sub_even_imag_entity_77ffaad0ab;

architecture structural of sub_even_imag_entity_77ffaad0ab is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x9: std_logic;
  signal clk_1_sg_x9: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x12: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(17 downto 0);

begin
  reinterpret1_output_port_net_x11 <= a;
  reinterpret1_output_port_net_x12 <= b;
  ce_1_sg_x9 <= ce_1;
  clk_1_sg_x9 <= clk_1;
  dout <= reinterpret1_output_port_net_x13;

  a_debus_e3ba56e22c: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret1_output_port_net_x11,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_18f6f1cec46d694e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x9,
      ce => ce_1_sg_x9,
      clk => clk_1_sg_x9,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  b_debus_0860deab4b: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret1_output_port_net_x12,
      msb_lsb_out1 => reinterpret1_output_port_net_x9
    );

  op_bussify_8134ef1c53: entity work.op_bussify_entity_a0c10d7209
    port map (
      in1 => addsub1_s_net_x0,
      bus_out => reinterpret1_output_port_net_x13
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/hilbert0"

entity hilbert0_entity_47cbdf1a3e is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    even: out std_logic_vector(35 downto 0); 
    odd: out std_logic_vector(35 downto 0)
  );
end hilbert0_entity_47cbdf1a3e;

architecture structural of hilbert0_entity_47cbdf1a3e is
  signal ce_1_sg_x11: std_logic;
  signal clk_1_sg_x11: std_logic;
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concat_y_net_x2: std_logic_vector(35 downto 0);
  signal concat_y_net_x3: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(75 downto 0);
  signal mux0_y_net_x1: std_logic_vector(35 downto 0);
  signal mux1_y_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x12: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);

begin
  mux0_y_net_x1 <= a;
  mux1_y_net_x1 <= b;
  ce_1_sg_x11 <= ce_1;
  clk_1_sg_x11 <= clk_1;
  even <= reinterpret_out_output_port_net_x5;
  odd <= reinterpret_out_output_port_net_x6;

  add_even_real_d02be0cdd9: entity work.add_even_real_entity_d02be0cdd9
    port map (
      a => reinterpret2_output_port_net_x6,
      b => reinterpret2_output_port_net_x7,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x3
    );

  add_odd_real_be4875c231: entity work.add_even_real_entity_d02be0cdd9
    port map (
      a => reinterpret1_output_port_net_x11,
      b => reinterpret1_output_port_net_x12,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x7
    );

  bus_convert_6fcb7792a1: entity work.bus_convert_entity_6fcb7792a1
    port map (
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      din => concatenate_y_net_x5,
      dout => concatenate_y_net_x4
    );

  bus_expand_26ad604baf: entity work.bus_expand_entity_26ad604baf
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

  bus_expand_a_e0cf78c6cc: entity work.bus_expand_a_entity_e0cf78c6cc
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => reinterpret2_output_port_net_x6
    );

  bus_expand_b_f861987b0d: entity work.bus_expand_a_entity_e0cf78c6cc
    port map (
      bus_in => reinterpret_out_output_port_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x12,
      msb_out2 => reinterpret2_output_port_net_x7
    );

  bus_scale_472dd14792: entity work.bus_scale_entity_472dd14792
    port map (
      din => concat_y_net_x1,
      dout => concatenate_y_net_x5
    );

  concat: entity work.concat_2aea51ccde
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net_x3,
      in1 => reinterpret1_output_port_net_x4,
      in2 => reinterpret1_output_port_net_x13,
      in3 => reinterpret1_output_port_net_x7,
      y => concat_y_net_x1
    );

  munge_a_40c03aaddb: entity work.munge_a_entity_40c03aaddb
    port map (
      din => mux0_y_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_b_a95bce3af9: entity work.munge_a_entity_40c03aaddb
    port map (
      din => mux1_y_net_x1,
      dout => reinterpret_out_output_port_net_x2
    );

  munge_even_c0db61d0d5: entity work.munge_a_entity_40c03aaddb
    port map (
      din => concat_y_net_x2,
      dout => reinterpret_out_output_port_net_x5
    );

  munge_odd_3740c036f1: entity work.munge_a_entity_40c03aaddb
    port map (
      din => concat_y_net_x3,
      dout => reinterpret_out_output_port_net_x6
    );

  ri_to_c1_e86063d3a1: entity work.ri_to_c_entity_2b066e56b4
    port map (
      im => reinterpret3_output_port_net_x1,
      re => reinterpret1_output_port_net_x1,
      c => concat_y_net_x3
    );

  ri_to_c_2b066e56b4: entity work.ri_to_c_entity_2b066e56b4
    port map (
      im => reinterpret2_output_port_net_x1,
      re => reinterpret4_output_port_net_x1,
      c => concat_y_net_x2
    );

  sub_even_imag_77ffaad0ab: entity work.sub_even_imag_entity_77ffaad0ab
    port map (
      a => reinterpret1_output_port_net_x11,
      b => reinterpret1_output_port_net_x12,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x13
    );

  sub_odd_imag_4941b0550d: entity work.sub_even_imag_entity_77ffaad0ab
    port map (
      a => reinterpret2_output_port_net_x7,
      b => reinterpret2_output_port_net_x6,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/mirror_spectrum/complex_conj0/imag_negate/bussify"

entity bussify_entity_427b04c969 is
  port (
    in1: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(17 downto 0)
  );
end bussify_entity_427b04c969;

architecture structural of bussify_entity_427b04c969 is
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);

begin
  neg1_op_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => neg1_op_net_x0,
      output_port => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/mirror_spectrum/complex_conj0/imag_negate"

entity imag_negate_entity_fb3ca9c1b2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(17 downto 0); 
    dout: out std_logic_vector(17 downto 0)
  );
end imag_negate_entity_fb3ca9c1b2;

architecture structural of imag_negate_entity_fb3ca9c1b2 is
  signal ce_1_sg_x22: std_logic;
  signal clk_1_sg_x22: std_logic;
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x22 <= ce_1;
  clk_1_sg_x22 <= clk_1;
  reinterpret1_output_port_net_x4 <= din;
  dout <= reinterpret1_output_port_net_x5;

  bussify_427b04c969: entity work.bussify_entity_427b04c969
    port map (
      in1 => neg1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x5
    );

  debus_c3e923df74: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret1_output_port_net_x4,
      msb_lsb_out1 => reinterpret1_output_port_net_x3
    );

  neg1: entity work.negate_f983e30a8b
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      ip => reinterpret1_output_port_net_x3,
      op => neg1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/mirror_spectrum/complex_conj0"

entity complex_conj0_entity_786e23abb9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    z: in std_logic_vector(35 downto 0); 
    z_x0: out std_logic_vector(35 downto 0)
  );
end complex_conj0_entity_786e23abb9;

architecture structural of complex_conj0_entity_786e23abb9 is
  signal ce_1_sg_x23: std_logic;
  signal clk_1_sg_x23: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal d3_q_net_x1: std_logic_vector(35 downto 0);
  signal real_delay_q_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x23 <= ce_1;
  clk_1_sg_x23 <= clk_1;
  d3_q_net_x1 <= z;
  z_x0 <= reinterpret_out_output_port_net_x2;

  bus_create_eb41049930: entity work.join_entity_dce4ac7e98
    port map (
      in1 => real_delay_q_net_x0,
      in2 => reinterpret1_output_port_net_x5,
      bus_out => concatenate_y_net_x2
    );

  bus_expand_379143f788: entity work.bus_expand_a_entity_e0cf78c6cc
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  imag_negate_fb3ca9c1b2: entity work.imag_negate_entity_fb3ca9c1b2
    port map (
      ce_1 => ce_1_sg_x23,
      clk_1 => clk_1_sg_x23,
      din => reinterpret1_output_port_net_x4,
      dout => reinterpret1_output_port_net_x5
    );

  munge_in_0f3d9693f0: entity work.munge_a_entity_40c03aaddb
    port map (
      din => d3_q_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_out_da2e9f6c3a: entity work.munge_a_entity_40c03aaddb
    port map (
      din => concatenate_y_net_x2,
      dout => reinterpret_out_output_port_net_x2
    );

  real_delay: entity work.delay_6699ee0916
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x0,
      q => real_delay_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/mirror_spectrum"

entity mirror_spectrum_entity_a832d647f2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    din1: in std_logic_vector(35 downto 0); 
    din2: in std_logic_vector(35 downto 0); 
    din3: in std_logic_vector(35 downto 0); 
    reo_in0: in std_logic_vector(35 downto 0); 
    reo_in1: in std_logic_vector(35 downto 0); 
    reo_in2: in std_logic_vector(35 downto 0); 
    reo_in3: in std_logic_vector(35 downto 0); 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    dout1: out std_logic_vector(35 downto 0); 
    dout2: out std_logic_vector(35 downto 0); 
    dout3: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end mirror_spectrum_entity_a832d647f2;

architecture structural of mirror_spectrum_entity_a832d647f2 is
  signal ce_1_sg_x30: std_logic;
  signal clk_1_sg_x30: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal d3_q_net_x2: std_logic_vector(35 downto 0);
  signal d4_q_net_x2: std_logic_vector(35 downto 0);
  signal d5_q_net_x2: std_logic_vector(35 downto 0);
  signal d6_q_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net: std_logic_vector(35 downto 0);
  signal delay1_q_net: std_logic_vector(35 downto 0);
  signal delay2_q_net: std_logic_vector(35 downto 0);
  signal delay3_q_net: std_logic_vector(35 downto 0);
  signal mux0_y_net_x0: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux2_y_net_x0: std_logic_vector(35 downto 0);
  signal mux3_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x0: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x9: std_logic_vector(35 downto 0);
  signal relational_op_net: std_logic;
  signal sync_delay0_q_net: std_logic;
  signal sync_delay1_q_net_x0: std_logic;

begin
  ce_1_sg_x30 <= ce_1;
  clk_1_sg_x30 <= clk_1;
  ram_data_out_net_x2 <= din0;
  ram_data_out_net_x3 <= din1;
  reinterpret_out_output_port_net_x9 <= din2;
  reinterpret_out_output_port_net_x10 <= din3;
  d3_q_net_x2 <= reo_in0;
  d4_q_net_x2 <= reo_in1;
  d5_q_net_x2 <= reo_in2;
  d6_q_net_x2 <= reo_in3;
  mux_y_net_x0 <= sync;
  dout0 <= mux0_y_net_x0;
  dout1 <= mux1_y_net_x0;
  dout2 <= mux2_y_net_x0;
  dout3 <= mux3_y_net_x0;
  sync_out <= sync_delay1_q_net_x0;

  complex_conj0_786e23abb9: entity work.complex_conj0_entity_786e23abb9
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      z => d3_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x2
    );

  complex_conj1_8286c9f2d5: entity work.complex_conj0_entity_786e23abb9
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      z => d4_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x6
    );

  complex_conj2_9f530b79ff: entity work.complex_conj0_entity_786e23abb9
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      z => d5_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x7
    );

  complex_conj3_94a422fdb8: entity work.complex_conj0_entity_786e23abb9
    port map (
      ce_1 => ce_1_sg_x30,
      clk_1 => clk_1_sg_x30,
      z => d6_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x8
    );

  constant_x0: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      en => "1",
      rst(0) => sync_delay0_q_net,
      op => counter_op_net
    );

  delay0: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d => ram_data_out_net_x2,
      q => delay0_q_net
    );

  delay1: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d => ram_data_out_net_x3,
      q => delay1_q_net
    );

  delay2: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d => reinterpret_out_output_port_net_x9,
      q => delay2_q_net
    );

  delay3: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d => reinterpret_out_output_port_net_x10,
      q => delay3_q_net
    );

  mux0: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d0 => delay0_q_net,
      d1 => reinterpret_out_output_port_net_x2,
      sel(0) => relational_op_net,
      y => mux0_y_net_x0
    );

  mux1: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d0 => delay1_q_net,
      d1 => reinterpret_out_output_port_net_x6,
      sel(0) => relational_op_net,
      y => mux1_y_net_x0
    );

  mux2: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d0 => delay2_q_net,
      d1 => reinterpret_out_output_port_net_x7,
      sel(0) => relational_op_net,
      y => mux2_y_net_x0
    );

  mux3: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d0 => delay3_q_net,
      d1 => reinterpret_out_output_port_net_x8,
      sel(0) => relational_op_net,
      y => mux3_y_net_x0
    );

  relational: entity work.relational_54e7975215
    port map (
      a => counter_op_net,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  sync_delay0: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => sync_delay0_q_net
    );

  sync_delay1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d(0) => sync_delay0_q_net,
      q(0) => sync_delay1_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/reorder_even/sync_delay_en"

entity sync_delay_en_entity_0faaba4daf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_en_entity_0faaba4daf;

architecture structural of sync_delay_en_entity_0faaba4daf is
  signal ce_1_sg_x31: std_logic;
  signal clk_1_sg_x31: std_logic;
  signal constant1_op_net: std_logic_vector(12 downto 0);
  signal constant2_op_net: std_logic_vector(12 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal logical1_y_net: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x0: std_logic;
  signal or_y_net_x0: std_logic;
  signal pre_sync_delay_q_net_x0: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x31 <= ce_1;
  clk_1_sg_x31 <= clk_1;
  or_y_net_x0 <= en;
  pre_sync_delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x0;

  constant1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_50be3b5040
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_461fd5d45cff2f9b",
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x31,
      clk => clk_1_sg_x31,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical1_y_net,
      load(0) => pre_sync_delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net,
      d1(0) => or_y_net_x0,
      y(0) => logical1_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x0
    );

  relational: entity work.relational_6dfa374756
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_2550da35d2
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/reorder_even"

entity reorder_even_entity_579a759212 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end reorder_even_entity_579a759212;

architecture structural of reorder_even_entity_579a759212 is
  signal bram0_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ce_1_sg_x32: std_logic;
  signal clk_1_sg_x32: std_logic;
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we_q_net: std_logic;
  signal en_even_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic;
  signal or_y_net_x0: std_logic;
  signal post_sync_delay_q_net_x0: std_logic;
  signal pre_sync_delay_q_net_x0: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x32 <= ce_1;
  clk_1_sg_x32 <= clk_1;
  reinterpret2_output_port_net_x0 <= din0;
  en_even_op_net_x0 <= en;
  delay0_q_net_x0 <= sync;
  dout0 <= bram0_data_out_net_x0;
  sync_out <= post_sync_delay_q_net_x0;

  bram0: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      data_in => delay_din0_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram0_data_out_net_x0
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 8191,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      count_limited => 0,
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      en(0) => en_even_op_net_x0,
      rst(0) => delay0_q_net_x0,
      op => counter_op_net
    );

  delay_d0: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      d => reinterpret2_output_port_net_x0,
      q => delay_din0_q_net
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_21355083c1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      d(0) => en_even_op_net_x0,
      q(0) => delay_we_q_net
    );

  map1: entity work.xlsprom_dist_fft_core
    generic map (
      addr_width => 12,
      c_address_width => 12,
      c_width => 12,
      core_name0 => "dmg_72_08915946f5ebdf9c",
      latency => 0
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      en => "1",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net
    );

  or_x0: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => delay_we_q_net,
      y(0) => or_y_net_x0
    );

  post_sync_delay: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => post_sync_delay_q_net_x0
    );

  pre_sync_delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      d(0) => delay0_q_net_x0,
      q(0) => pre_sync_delay_q_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

  sync_delay_en_0faaba4daf: entity work.sync_delay_en_entity_0faaba4daf
    port map (
      ce_1 => ce_1_sg_x32,
      clk_1 => clk_1_sg_x32,
      en => or_y_net_x0,
      in_x0 => pre_sync_delay_q_net_x0,
      out_x0 => mux_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/reorder_odd"

entity reorder_odd_entity_a1b8b27aff is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0)
  );
end reorder_odd_entity_a1b8b27aff;

architecture structural of reorder_odd_entity_a1b8b27aff is
  signal bram0_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ce_1_sg_x33: std_logic;
  signal clk_1_sg_x33: std_logic;
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we_q_net: std_logic;
  signal en_odd_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x33 <= ce_1;
  clk_1_sg_x33 <= clk_1;
  reinterpret1_output_port_net_x0 <= din0;
  en_odd_op_net_x0 <= en;
  delay0_q_net_x1 <= sync;
  dout0 <= bram0_data_out_net_x0;

  bram0: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      data_in => delay_din0_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram0_data_out_net_x0
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 8191,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      count_limited => 0,
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      clr => '0',
      en(0) => en_odd_op_net_x0,
      rst(0) => delay0_q_net_x1,
      op => counter_op_net
    );

  delay_d0: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => delay_din0_q_net
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_21355083c1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      clr => '0',
      d(0) => en_odd_op_net_x0,
      q(0) => delay_we_q_net
    );

  map1: entity work.xlsprom_dist_fft_core
    generic map (
      addr_width => 12,
      c_address_width => 12,
      c_width => 12,
      core_name0 => "dmg_72_b5cea772b1c370b5",
      latency => 0
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      en => "1",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/reorder_out"

entity reorder_out_entity_9cf6a341de is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    din1: in std_logic_vector(35 downto 0); 
    din2: in std_logic_vector(35 downto 0); 
    din3: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    dout1: out std_logic_vector(35 downto 0); 
    dout2: out std_logic_vector(35 downto 0); 
    dout3: out std_logic_vector(35 downto 0)
  );
end reorder_out_entity_9cf6a341de;

architecture structural of reorder_out_entity_9cf6a341de is
  signal bram0_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ce_1_sg_x34: std_logic;
  signal clk_1_sg_x34: std_logic;
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net: std_logic_vector(35 downto 0);
  signal delay_din1_q_net: std_logic_vector(35 downto 0);
  signal delay_din2_q_net: std_logic_vector(35 downto 0);
  signal delay_din3_q_net: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we_q_net: std_logic;
  signal en_out_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal mux_y_net_x1: std_logic;
  signal ram_data_out_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x12: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x34 <= ce_1;
  clk_1_sg_x34 <= clk_1;
  ram_data_out_net_x4 <= din0;
  ram_data_out_net_x5 <= din1;
  reinterpret_out_output_port_net_x11 <= din2;
  reinterpret_out_output_port_net_x12 <= din3;
  en_out_op_net_x0 <= en;
  mux_y_net_x1 <= sync;
  dout0 <= bram0_data_out_net_x0;
  dout1 <= bram1_data_out_net_x0;
  dout2 <= bram2_data_out_net_x0;
  dout3 <= bram3_data_out_net_x0;

  bram0: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      data_in => delay_din0_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram0_data_out_net_x0
    );

  bram1: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      data_in => delay_din1_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram1_data_out_net_x0
    );

  bram2: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      data_in => delay_din2_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram2_data_out_net_x0
    );

  bram3: entity work.xlspram_fft_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_f0e087429b44571a",
      latency => 2
    )
    port map (
      addr => mux_y_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      data_in => delay_din3_q_net,
      en => "1",
      rst => "0",
      we(0) => delay_we_q_net,
      data_out => bram3_data_out_net_x0
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 8191,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      count_limited => 0,
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      en(0) => en_out_op_net_x0,
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  delay_d0: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => ram_data_out_net_x4,
      q => delay_din0_q_net
    );

  delay_din1: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => ram_data_out_net_x5,
      q => delay_din1_q_net
    );

  delay_din2: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => reinterpret_out_output_port_net_x11,
      q => delay_din2_q_net
    );

  delay_din3: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => reinterpret_out_output_port_net_x12,
      q => delay_din3_q_net
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_21355083c1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d(0) => en_out_op_net_x0,
      q(0) => delay_we_q_net
    );

  map1: entity work.xlsprom_dist_fft_core
    generic map (
      addr_width => 12,
      c_address_width => 12,
      c_width => 12,
      core_name0 => "dmg_72_f54beabec7472b25",
      latency => 0
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      en => "1",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x/sync_delay"

entity sync_delay_entity_a3385278ea is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_a3385278ea;

architecture structural of sync_delay_entity_a3385278ea is
  signal ce_1_sg_x35: std_logic;
  signal clk_1_sg_x35: std_logic;
  signal constant1_op_net: std_logic_vector(12 downto 0);
  signal constant2_op_net: std_logic_vector(12 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal d2_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x2: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x35 <= ce_1;
  clk_1_sg_x35 <= clk_1;
  d2_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x2;

  constant1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_50be3b5040
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_461fd5d45cff2f9b",
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => d2_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => d2_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => d2_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x2
    );

  relational: entity work.relational_6dfa374756
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_2550da35d2
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/bi_real_unscr_4x"

entity bi_real_unscr_4x_entity_8d809182bf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    even: in std_logic_vector(35 downto 0); 
    odd: in std_logic_vector(35 downto 0); 
    sync: in std_logic; 
    pol1_out: out std_logic_vector(35 downto 0); 
    pol2_out: out std_logic_vector(35 downto 0); 
    pol3_out: out std_logic_vector(35 downto 0); 
    pol4_out: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end bi_real_unscr_4x_entity_8d809182bf;

architecture structural of bi_real_unscr_4x_entity_8d809182bf is
  signal bram0_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram0_data_out_net_x1: std_logic_vector(35 downto 0);
  signal bram0_data_out_net_x2: std_logic_vector(35 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(35 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(35 downto 0);
  signal c0_op_net: std_logic_vector(12 downto 0);
  signal c1_op_net: std_logic_vector(12 downto 0);
  signal ce_1_sg_x36: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal count_op_net: std_logic_vector(12 downto 0);
  signal d0_q_net: std_logic_vector(35 downto 0);
  signal d2_q_net_x0: std_logic;
  signal d3_q_net_x2: std_logic_vector(35 downto 0);
  signal d4_q_net_x2: std_logic_vector(35 downto 0);
  signal d5_q_net_x2: std_logic_vector(35 downto 0);
  signal d6_q_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal en_even_op_net_x0: std_logic;
  signal en_odd_op_net_x0: std_logic;
  signal en_out_op_net_x0: std_logic;
  signal mux0_y_net_x1: std_logic_vector(35 downto 0);
  signal mux0_y_net_x2: std_logic_vector(35 downto 0);
  signal mux1_y_net_x1: std_logic_vector(35 downto 0);
  signal mux1_y_net_x2: std_logic_vector(35 downto 0);
  signal mux2_y_net_x1: std_logic_vector(35 downto 0);
  signal mux2_y_net_x2: std_logic_vector(35 downto 0);
  signal mux3_y_net_x1: std_logic_vector(35 downto 0);
  signal mux3_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal post_sync_delay_q_net_x0: std_logic;
  signal r0_op_net: std_logic;
  signal r1_op_net: std_logic;
  signal ram_data_out_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);
  signal sync_delay1_q_net_x1: std_logic;

begin
  ce_1_sg_x36 <= ce_1;
  clk_1_sg_x36 <= clk_1;
  reinterpret2_output_port_net_x1 <= even;
  reinterpret1_output_port_net_x1 <= odd;
  delay0_q_net_x2 <= sync;
  pol1_out <= mux0_y_net_x2;
  pol2_out <= mux1_y_net_x2;
  pol3_out <= mux2_y_net_x2;
  pol4_out <= mux3_y_net_x2;
  sync_out <= sync_delay1_q_net_x1;

  c0: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => c0_op_net
    );

  c1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => c1_op_net
    );

  count: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      en => "1",
      rst(0) => post_sync_delay_q_net_x0,
      op => count_op_net
    );

  d0: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d => bram0_data_out_net_x1,
      q => d0_q_net
    );

  d2: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d(0) => post_sync_delay_q_net_x0,
      q(0) => d2_q_net_x0
    );

  d3: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d => bram0_data_out_net_x2,
      q => d3_q_net_x2
    );

  d4: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d => bram1_data_out_net_x0,
      q => d4_q_net_x2
    );

  d5: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d => bram2_data_out_net_x0,
      q => d5_q_net_x2
    );

  d6: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d => bram3_data_out_net_x0,
      q => d6_q_net_x2
    );

  delay0_4675455b89: entity work.delay0_entity_4675455b89
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din => reinterpret_out_output_port_net_x5,
      dout => ram_data_out_net_x4
    );

  delay1_4221f778ec: entity work.delay0_entity_4675455b89
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din => reinterpret_out_output_port_net_x6,
      dout => ram_data_out_net_x5
    );

  en_even: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_even_op_net_x0
    );

  en_odd: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_odd_op_net_x0
    );

  en_out: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_out_op_net_x0
    );

  hilbert0_47cbdf1a3e: entity work.hilbert0_entity_47cbdf1a3e
    port map (
      a => mux0_y_net_x1,
      b => mux1_y_net_x1,
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      even => reinterpret_out_output_port_net_x5,
      odd => reinterpret_out_output_port_net_x6
    );

  hilbert1_9f3ab3bb55: entity work.hilbert0_entity_47cbdf1a3e
    port map (
      a => mux2_y_net_x1,
      b => mux3_y_net_x1,
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      even => reinterpret_out_output_port_net_x11,
      odd => reinterpret_out_output_port_net_x12
    );

  mirror_spectrum_a832d647f2: entity work.mirror_spectrum_entity_a832d647f2
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din0 => ram_data_out_net_x4,
      din1 => ram_data_out_net_x5,
      din2 => reinterpret_out_output_port_net_x11,
      din3 => reinterpret_out_output_port_net_x12,
      reo_in0 => d3_q_net_x2,
      reo_in1 => d4_q_net_x2,
      reo_in2 => d5_q_net_x2,
      reo_in3 => d6_q_net_x2,
      sync => mux_y_net_x2,
      dout0 => mux0_y_net_x2,
      dout1 => mux1_y_net_x2,
      dout2 => mux2_y_net_x2,
      dout3 => mux3_y_net_x2,
      sync_out => sync_delay1_q_net_x1
    );

  mux0: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d0 => bram0_data_out_net_x0,
      d1 => d0_q_net,
      sel(0) => r0_op_net,
      y => mux0_y_net_x1
    );

  mux1: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d0 => d0_q_net,
      d1 => bram0_data_out_net_x0,
      sel(0) => r1_op_net,
      y => mux1_y_net_x1
    );

  mux2: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d0 => bram0_data_out_net_x0,
      d1 => d0_q_net,
      sel(0) => r1_op_net,
      y => mux2_y_net_x1
    );

  mux3: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      d0 => d0_q_net,
      d1 => bram0_data_out_net_x0,
      sel(0) => r0_op_net,
      y => mux3_y_net_x1
    );

  r0: entity work.relational_6dfa374756
    port map (
      a => c0_op_net,
      b => count_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => r0_op_net
    );

  r1: entity work.relational_6dfa374756
    port map (
      a => count_op_net,
      b => c1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => r1_op_net
    );

  reorder_even_579a759212: entity work.reorder_even_entity_579a759212
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din0 => reinterpret2_output_port_net_x1,
      en => en_even_op_net_x0,
      sync => delay0_q_net_x2,
      dout0 => bram0_data_out_net_x0,
      sync_out => post_sync_delay_q_net_x0
    );

  reorder_odd_a1b8b27aff: entity work.reorder_odd_entity_a1b8b27aff
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din0 => reinterpret1_output_port_net_x1,
      en => en_odd_op_net_x0,
      sync => delay0_q_net_x2,
      dout0 => bram0_data_out_net_x1
    );

  reorder_out_9cf6a341de: entity work.reorder_out_entity_9cf6a341de
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      din0 => ram_data_out_net_x4,
      din1 => ram_data_out_net_x5,
      din2 => reinterpret_out_output_port_net_x11,
      din3 => reinterpret_out_output_port_net_x12,
      en => en_out_op_net_x0,
      sync => mux_y_net_x2,
      dout0 => bram0_data_out_net_x2,
      dout1 => bram1_data_out_net_x0,
      dout2 => bram2_data_out_net_x0,
      dout3 => bram3_data_out_net_x0
    );

  sync_delay_a3385278ea: entity work.sync_delay_entity_a3385278ea
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      in_x0 => d2_q_net_x0,
      out_x0 => mux_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_add/a_debus"

entity a_debus_entity_c0242f8ce0 is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out2: out std_logic_vector(17 downto 0)
  );
end a_debus_entity_c0242f8ce0;

architecture structural of a_debus_entity_c0242f8ce0 is
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);

begin
  ram_data_out_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => ram_data_out_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => ram_data_out_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_add/op_bussify"

entity op_bussify_entity_8ee3422350 is
  port (
    in1: in std_logic_vector(18 downto 0); 
    in2: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(37 downto 0)
  );
end op_bussify_entity_8ee3422350;

architecture structural of op_bussify_entity_8ee3422350 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(37 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(18 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  addsub2_s_net_x0 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_5a12f8f9be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub2_s_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_add"

entity bus_add_entity_695cb26b69 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(37 downto 0)
  );
end bus_add_entity_695cb26b69;

architecture structural of bus_add_entity_695cb26b69 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x37: std_logic;
  signal clk_1_sg_x37: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(37 downto 0);
  signal mux_y_net_x1: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  ram_data_out_net_x1 <= a;
  mux_y_net_x1 <= b;
  ce_1_sg_x37 <= ce_1;
  clk_1_sg_x37 <= clk_1;
  dout <= concatenate_y_net_x1;

  a_debus_c0242f8ce0: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => ram_data_out_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_0b9daa5d24360c6e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_0b9daa5d24360c6e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_3efe4bc196: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => mux_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_8ee3422350: entity work.op_bussify_entity_8ee3422350
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_convert/conv1/convert"

entity convert_entity_1c9b149e9c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(19 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end convert_entity_1c9b149e9c;

architecture structural of convert_entity_1c9b149e9c is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x38: std_logic;
  signal clk_1_sg_x38: std_logic;
  signal concat_y_net: std_logic_vector(20 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(20 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(19 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x38 <= ce_1;
  clk_1_sg_x38 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.addsub_b96bfee539
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x38,
      clk => clk_1_sg_x38,
      clr => '0',
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 19,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_c615d93998
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_convert/conv1"

entity conv1_entity_32aefab339 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(19 downto 0); 
    dout: out std_logic_vector(17 downto 0); 
    of_x0: out std_logic
  );
end conv1_entity_32aefab339;

architecture structural of conv1_entity_32aefab339 is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal all_0s_y_net: std_logic;
  signal all_1s_y_net: std_logic;
  signal and_y_net_x0: std_logic;
  signal ce_1_sg_x39: std_logic;
  signal clk_1_sg_x39: std_logic;
  signal invert1_op_net: std_logic;
  signal invert2_op_net: std_logic;
  signal reinterpret4_output_port_net_x1: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic;

begin
  ce_1_sg_x39 <= ce_1;
  clk_1_sg_x39 <= clk_1;
  reinterpret4_output_port_net_x1 <= din;
  dout <= adder_s_net_x5;
  of_x0 <= and_y_net_x0;

  all_0s: entity work.logical_5bc1b3bb27
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d0(0) => invert1_op_net,
      d1(0) => invert2_op_net,
      y(0) => all_0s_y_net
    );

  all_1s: entity work.logical_5bc1b3bb27
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d0(0) => slice1_y_net,
      d1(0) => slice2_y_net,
      y(0) => all_1s_y_net
    );

  and_x0: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => all_0s_y_net,
      d1(0) => all_1s_y_net,
      y(0) => and_y_net_x0
    );

  convert_1c9b149e9c: entity work.convert_entity_1c9b149e9c
    port map (
      ce_1 => ce_1_sg_x39,
      clk_1 => clk_1_sg_x39,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  invert1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      ip(0) => slice1_y_net,
      op(0) => invert1_op_net
    );

  invert2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      ip(0) => slice2_y_net,
      op(0) => invert2_op_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 19,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 18,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_convert/debus"

entity debus_entity_71deb38b98 is
  port (
    bus_in: in std_logic_vector(79 downto 0); 
    lsb_out1: out std_logic_vector(19 downto 0); 
    msb_out4: out std_logic_vector(19 downto 0); 
    out2: out std_logic_vector(19 downto 0); 
    out3: out std_logic_vector(19 downto 0)
  );
end debus_entity_71deb38b98;

architecture structural of debus_entity_71deb38b98 is
  signal mux_y_net_x0: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic_vector(19 downto 0);
  signal slice2_y_net: std_logic_vector(19 downto 0);
  signal slice3_y_net: std_logic_vector(19 downto 0);
  signal slice4_y_net: std_logic_vector(19 downto 0);

begin
  mux_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out4 <= reinterpret4_output_port_net_x2;
  out2 <= reinterpret2_output_port_net_x2;
  out3 <= reinterpret3_output_port_net_x2;

  reinterpret1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  reinterpret3: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x2
    );

  reinterpret4: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 19,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => mux_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 39,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => mux_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 59,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => mux_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 79,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => mux_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_convert/of_bussify"

entity of_bussify_entity_be16087e66 is
  port (
    in1: in std_logic; 
    in2: in std_logic; 
    in3: in std_logic; 
    in4: in std_logic; 
    bus_out: out std_logic_vector(3 downto 0)
  );
end of_bussify_entity_be16087e66;

architecture structural of of_bussify_entity_be16087e66 is
  signal and_y_net_x4: std_logic;
  signal and_y_net_x5: std_logic;
  signal and_y_net_x6: std_logic;
  signal and_y_net_x7: std_logic;
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net: std_logic;
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic;
  signal reinterpret4_output_port_net: std_logic;

begin
  and_y_net_x4 <= in1;
  and_y_net_x5 <= in2;
  and_y_net_x6 <= in3;
  and_y_net_x7 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2(0) => reinterpret3_output_port_net,
      in3(0) => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => and_y_net_x4,
      output_port(0) => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => and_y_net_x5,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => and_y_net_x6,
      output_port(0) => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => and_y_net_x7,
      output_port(0) => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_convert"

entity bus_convert_entity_82369b5cdf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(71 downto 0); 
    overflow: out std_logic_vector(3 downto 0)
  );
end bus_convert_entity_82369b5cdf;

architecture structural of bus_convert_entity_82369b5cdf is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal adder_s_net_x8: std_logic_vector(17 downto 0);
  signal and_y_net_x4: std_logic;
  signal and_y_net_x5: std_logic;
  signal and_y_net_x6: std_logic;
  signal and_y_net_x7: std_logic;
  signal ce_1_sg_x46: std_logic;
  signal clk_1_sg_x46: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(3 downto 0);
  signal mux_y_net_x1: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x46 <= ce_1;
  clk_1_sg_x46 <= clk_1;
  mux_y_net_x1 <= din;
  dout <= concatenate_y_net_x2;
  overflow <= concatenate_y_net_x3;

  bussify_08dd535688: entity work.bussify_entity_1d06622102
    port map (
      in1 => adder_s_net_x5,
      in2 => adder_s_net_x6,
      in3 => adder_s_net_x7,
      in4 => adder_s_net_x8,
      bus_out => concatenate_y_net_x2
    );

  conv1_32aefab339: entity work.conv1_entity_32aefab339
    port map (
      ce_1 => ce_1_sg_x46,
      clk_1 => clk_1_sg_x46,
      din => reinterpret4_output_port_net_x2,
      dout => adder_s_net_x5,
      of_x0 => and_y_net_x4
    );

  conv2_449a6556a1: entity work.conv1_entity_32aefab339
    port map (
      ce_1 => ce_1_sg_x46,
      clk_1 => clk_1_sg_x46,
      din => reinterpret3_output_port_net_x2,
      dout => adder_s_net_x6,
      of_x0 => and_y_net_x5
    );

  conv3_fa7836b597: entity work.conv1_entity_32aefab339
    port map (
      ce_1 => ce_1_sg_x46,
      clk_1 => clk_1_sg_x46,
      din => reinterpret2_output_port_net_x2,
      dout => adder_s_net_x7,
      of_x0 => and_y_net_x6
    );

  conv4_6ba04c258a: entity work.conv1_entity_32aefab339
    port map (
      ce_1 => ce_1_sg_x46,
      clk_1 => clk_1_sg_x46,
      din => reinterpret1_output_port_net_x2,
      dout => adder_s_net_x8,
      of_x0 => and_y_net_x7
    );

  debus_71deb38b98: entity work.debus_entity_71deb38b98
    port map (
      bus_in => mux_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

  of_bussify_be16087e66: entity work.of_bussify_entity_be16087e66
    port map (
      in1 => and_y_net_x4,
      in2 => and_y_net_x5,
      in3 => and_y_net_x6,
      in4 => and_y_net_x7,
      bus_out => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_expand"

entity bus_expand_entity_2ff4545d65 is
  port (
    bus_in: in std_logic_vector(71 downto 0); 
    lsb_out1: out std_logic_vector(35 downto 0); 
    msb_out2: out std_logic_vector(35 downto 0)
  );
end bus_expand_entity_2ff4545d65;

architecture structural of bus_expand_entity_2ff4545d65 is
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);
  signal slice2_y_net: std_logic_vector(35 downto 0);

begin
  concatenate_y_net_x3 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 72,
      y_width => 36
    )
    port map (
      x => concatenate_y_net_x3,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 71,
      x_width => 72,
      y_width => 36
    )
    port map (
      x => concatenate_y_net_x3,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_norm0/bussify"

entity bussify_entity_6546069b97 is
  port (
    in1: in std_logic_vector(19 downto 0); 
    in2: in std_logic_vector(19 downto 0); 
    in3: in std_logic_vector(19 downto 0); 
    in4: in std_logic_vector(19 downto 0); 
    bus_out: out std_logic_vector(79 downto 0)
  );
end bussify_entity_6546069b97;

architecture structural of bussify_entity_6546069b97 is
  signal concatenate_y_net_x0: std_logic_vector(79 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(19 downto 0);

begin
  conv1_dout_net_x0 <= in1;
  conv2_dout_net_x0 <= in2;
  conv3_dout_net_x0 <= in3;
  conv4_dout_net_x0 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_f86ebb6084
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv1_dout_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv2_dout_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv3_dout_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv4_dout_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_norm0"

entity bus_norm0_entity_f70daa5f43 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_norm0_entity_f70daa5f43;

architecture structural of bus_norm0_entity_f70daa5f43 is
  signal ce_1_sg_x47: std_logic;
  signal clk_1_sg_x47: std_logic;
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(79 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x47 <= ce_1;
  clk_1_sg_x47 <= clk_1;
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x1;

  bussify_6546069b97: entity work.bussify_entity_6546069b97
    port map (
      in1 => conv1_dout_net_x0,
      in2 => conv2_dout_net_x0,
      in3 => conv3_dout_net_x0,
      in4 => conv4_dout_net_x0,
      bus_out => concatenate_y_net_x1
    );

  conv1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      din => reinterpret4_output_port_net_x0,
      en => "1",
      dout => conv1_dout_net_x0
    );

  conv2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      din => reinterpret3_output_port_net_x0,
      en => "1",
      dout => conv2_dout_net_x0
    );

  conv3: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      din => reinterpret2_output_port_net_x0,
      en => "1",
      dout => conv3_dout_net_x0
    );

  conv4: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      din => reinterpret1_output_port_net_x0,
      en => "1",
      dout => conv4_dout_net_x0
    );

  debus_81ba5a08bf: entity work.debus_entity_8ef01a3c6c
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_norm1/conv1"

entity conv1_entity_68a3012b52 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(18 downto 0); 
    out_x0: out std_logic_vector(19 downto 0)
  );
end conv1_entity_68a3012b52;

architecture structural of conv1_entity_68a3012b52 is
  signal adder_s_net_x4: std_logic_vector(19 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x48: std_logic;
  signal clk_1_sg_x48: std_logic;
  signal concat_y_net: std_logic_vector(19 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(19 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(18 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x48 <= ce_1;
  clk_1_sg_x48 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.addsub_ba2df6ec2d
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      clr => '0',
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_b366689086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 19,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_504cae28bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_b1e9d7c303
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_norm1"

entity bus_norm1_entity_1de1ca87af is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_norm1_entity_1de1ca87af;

architecture structural of bus_norm1_entity_1de1ca87af is
  signal adder_s_net_x4: std_logic_vector(19 downto 0);
  signal adder_s_net_x5: std_logic_vector(19 downto 0);
  signal adder_s_net_x6: std_logic_vector(19 downto 0);
  signal adder_s_net_x7: std_logic_vector(19 downto 0);
  signal ce_1_sg_x52: std_logic;
  signal clk_1_sg_x52: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x52 <= ce_1;
  clk_1_sg_x52 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_4efdd54be1: entity work.bussify_entity_6546069b97
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_68a3012b52: entity work.conv1_entity_68a3012b52
    port map (
      ce_1 => ce_1_sg_x52,
      clk_1 => clk_1_sg_x52,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_996d8a099f: entity work.conv1_entity_68a3012b52
    port map (
      ce_1 => ce_1_sg_x52,
      clk_1 => clk_1_sg_x52,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_2ae1d2527a: entity work.conv1_entity_68a3012b52
    port map (
      ce_1 => ce_1_sg_x52,
      clk_1 => clk_1_sg_x52,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_39eba9037a: entity work.conv1_entity_68a3012b52
    port map (
      ce_1 => ce_1_sg_x52,
      clk_1 => clk_1_sg_x52,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_422a9e88b5: entity work.debus_entity_3f078924c3
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_relational/a_debus"

entity a_debus_entity_45cbe64c62 is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    msb_lsb_out1: out std_logic_vector(3 downto 0)
  );
end a_debus_entity_45cbe64c62;

architecture structural of a_debus_entity_45cbe64c62 is
  signal constant_op_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net: std_logic_vector(3 downto 0);

begin
  constant_op_net_x0 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 4,
      y_width => 4
    )
    port map (
      x => constant_op_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_relational/bussify"

entity bussify_entity_a249a45e4d is
  port (
    in1: in std_logic; 
    bus_out: out std_logic
  );
end bussify_entity_a249a45e4d;

architecture structural of bussify_entity_a249a45e4d is
  signal reinterpret1_output_port_net_x0: std_logic;
  signal relational1_op_net_x0: std_logic;

begin
  relational1_op_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => relational1_op_net_x0,
      output_port(0) => reinterpret1_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_relational"

entity bus_relational_entity_53f1d0be84 is
  port (
    a: in std_logic_vector(3 downto 0); 
    b: in std_logic_vector(3 downto 0); 
    a_b: out std_logic
  );
end bus_relational_entity_53f1d0be84;

architecture structural of bus_relational_entity_53f1d0be84 is
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic;
  signal reinterpret_out_output_port_net_x1: std_logic_vector(3 downto 0);
  signal relational1_op_net_x0: std_logic;

begin
  constant_op_net_x1 <= a;
  reinterpret_out_output_port_net_x1 <= b;
  a_b <= reinterpret1_output_port_net_x3;

  a_debus_45cbe64c62: entity work.a_debus_entity_45cbe64c62
    port map (
      bus_in => constant_op_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  b_debus_cedd82b2f6: entity work.a_debus_entity_45cbe64c62
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  bussify_a249a45e4d: entity work.bussify_entity_a249a45e4d
    port map (
      in1 => relational1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x3
    );

  relational1: entity work.relational_d930162434
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/bus_sub"

entity bus_sub_entity_2925aed405 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(37 downto 0)
  );
end bus_sub_entity_2925aed405;

architecture structural of bus_sub_entity_2925aed405 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x53: std_logic;
  signal clk_1_sg_x53: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(37 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  ram_data_out_net_x3 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x53 <= ce_1;
  clk_1_sg_x53 <= clk_1;
  dout <= concatenate_y_net_x1;

  a_debus_eaae6ef99a: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => ram_data_out_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_c9b173d075a3b6d7",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_c9b173d075a3b6d7",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_5cd917c1e7: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => mux_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_a5fdf8aaa8: entity work.op_bussify_entity_8ee3422350
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/munge/join"

entity join_entity_23d6dd178e is
  port (
    in1: in std_logic_vector(1 downto 0); 
    in2: in std_logic_vector(1 downto 0); 
    bus_out: out std_logic_vector(3 downto 0)
  );
end join_entity_23d6dd178e;

architecture structural of join_entity_23d6dd178e is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(1 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(1 downto 0);

begin
  reinterpret2_output_port_net_x1 <= in1;
  reinterpret1_output_port_net_x1 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret1_output_port_net_x1,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/munge/split"

entity split_entity_3865d2d8ca is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    lsb_out1: out std_logic_vector(1 downto 0); 
    msb_out2: out std_logic_vector(1 downto 0)
  );
end split_entity_3865d2d8ca;

architecture structural of split_entity_3865d2d8ca is
  signal reinterpret1_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net: std_logic_vector(1 downto 0);
  signal slice2_y_net: std_logic_vector(1 downto 0);

begin
  reinterpret_output_port_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out2 <= reinterpret2_output_port_net_x2;

  reinterpret1: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => reinterpret_output_port_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => reinterpret_output_port_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct/munge"

entity munge_entity_597456506f is
  port (
    din: in std_logic_vector(3 downto 0); 
    dout: out std_logic_vector(3 downto 0)
  );
end munge_entity_597456506f;

architecture structural of munge_entity_597456506f is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(3 downto 0);

begin
  concatenate_y_net_x4 <= din;
  dout <= reinterpret_out_output_port_net_x2;

  join_23d6dd178e: entity work.join_entity_23d6dd178e
    port map (
      in1 => reinterpret2_output_port_net_x2,
      in2 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x0
    );

  reinterpret: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x4,
      output_port => reinterpret_output_port_net_x0
    );

  reinterpret_out: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x0,
      output_port => reinterpret_out_output_port_net_x2
    );

  split_3865d2d8ca: entity work.split_entity_3865d2d8ca
    port map (
      bus_in => reinterpret_output_port_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1/butterfly_direct"

entity butterfly_direct_entity_4d29c42dd2 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_4d29c42dd2;

architecture structural of butterfly_direct_entity_4d29c42dd2 is
  signal ce_1_sg_x54: std_logic;
  signal clk_1_sg_x54: std_logic;
  signal concat_y_net_x3: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x0: std_logic;
  signal mux_y_net_x1: std_logic_vector(79 downto 0);
  signal mux_y_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x4 <= a;
  mux_y_net_x4 <= b;
  ce_1_sg_x54 <= ce_1;
  clk_1_sg_x54 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x0 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x5;
  sync_out <= delay0_q_net_x0;

  bus_add_695cb26b69: entity work.bus_add_entity_695cb26b69
    port map (
      a => ram_data_out_net_x4,
      b => mux_y_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      dout => concatenate_y_net_x1
    );

  bus_convert_82369b5cdf: entity work.bus_convert_entity_82369b5cdf
    port map (
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x3,
      overflow => concatenate_y_net_x4
    );

  bus_expand_2ff4545d65: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_f70daa5f43: entity work.bus_norm0_entity_f70daa5f43
    port map (
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x5
    );

  bus_norm1_1de1ca87af: entity work.bus_norm1_entity_1de1ca87af
    port map (
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_53f1d0be84: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x5
    );

  bus_scale_b2fbb42967: entity work.bus_scale_entity_472dd14792
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_2925aed405: entity work.bus_sub_entity_2925aed405
    port map (
      a => ram_data_out_net_x4,
      b => mux_y_net_x4,
      ce_1 => ce_1_sg_x54,
      clk_1 => clk_1_sg_x54,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_4822199898
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x1,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_597456506f: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x4,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_9ff8aec2dc
    port map (
      ce => ce_1_sg_x54,
      clk => clk_1_sg_x54,
      clr => '0',
      d0 => concatenate_y_net_x5,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_1"

entity fft_stage_1_entity_a0aa893753 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_1_entity_a0aa893753;

architecture structural of fft_stage_1_entity_a0aa893753 is
  signal ce_1_sg_x58: std_logic;
  signal clk_1_sg_x58: std_logic;
  signal constant_op_net_x0: std_logic;
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x0: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;
  signal sync_net_x0: std_logic;

begin
  ce_1_sg_x58 <= ce_1;
  clk_1_sg_x58 <= clk_1;
  reinterpret1_output_port_net_x1 <= in1;
  reinterpret1_output_port_net_x2 <= in2;
  constant_op_net_x0 <= of_in;
  fft_shift_net_x0 <= shift;
  sync_net_x0 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_4d29c42dd2: entity work.butterfly_direct_entity_4d29c42dd2
    port map (
      a => ram_data_out_net_x5,
      b => mux_y_net_x4,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x1,
      a_bw => reinterpret1_output_port_net_x6,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x5,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_125dc8e6a3ba8cad",
      op_arith => xlUnsigned,
      op_width => 13
    )
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      en => "1",
      rst(0) => sync_net_x0,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d(0) => sync_net_x0,
      q(0) => delay_q_net_x0
    );

  delay_b_307d66479a: entity work.delay0_entity_4675455b89
    port map (
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x5
    );

  delay_f_0b713717ed: entity work.delay0_entity_4675455b89
    port map (
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => reinterpret1_output_port_net_x2,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x5,
      d1(0) => constant_op_net_x0,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret1_output_port_net_x1,
      sel(0) => slice1_y_net,
      y => mux_y_net_x4
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d0 => reinterpret1_output_port_net_x1,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x0,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_6498f6a73b: entity work.sync_delay_entity_a3385278ea
    port map (
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_add/b_debus"

entity b_debus_entity_98717e8269 is
  port (
    bus_in: in std_logic_vector(37 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out2: out std_logic_vector(18 downto 0)
  );
end b_debus_entity_98717e8269;

architecture structural of b_debus_entity_98717e8269 is
  signal concatenate_y_net_x0: std_logic_vector(37 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 38,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 38,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_add/op_bussify"

entity op_bussify_entity_f21ce432ef is
  port (
    in1: in std_logic_vector(19 downto 0); 
    in2: in std_logic_vector(19 downto 0); 
    bus_out: out std_logic_vector(39 downto 0)
  );
end op_bussify_entity_f21ce432ef;

architecture structural of op_bussify_entity_f21ce432ef is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(19 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  addsub2_s_net_x0 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_9e724c4b50
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub2_s_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_add"

entity bus_add_entity_fda2dbc1e4 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(37 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(39 downto 0)
  );
end bus_add_entity_fda2dbc1e4;

architecture structural of bus_add_entity_fda2dbc1e4 is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal ce_1_sg_x59: std_logic;
  signal clk_1_sg_x59: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  reinterpret1_output_port_net_x3 <= a;
  concatenate_y_net_x2 <= b;
  ce_1_sg_x59 <= ce_1;
  clk_1_sg_x59 <= clk_1;
  dout <= concatenate_y_net_x3;

  a_debus_959fc4f209: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_6bbb8fb0d8f20abe",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_6bbb8fb0d8f20abe",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret1_output_port_net_x2,
      b => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_98717e8269: entity work.b_debus_entity_98717e8269
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_f21ce432ef: entity work.op_bussify_entity_f21ce432ef
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_convert/conv1/convert"

entity convert_entity_f7847c8c42 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(20 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end convert_entity_f7847c8c42;

architecture structural of convert_entity_f7847c8c42 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x60: std_logic;
  signal clk_1_sg_x60: std_logic;
  signal concat_y_net: std_logic_vector(21 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(21 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(20 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x60 <= ce_1;
  clk_1_sg_x60 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.addsub_6358c585f1
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 20,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_e6bc20c81b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_c84451c80b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_convert/conv1"

entity conv1_entity_11637058ac is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(20 downto 0); 
    dout: out std_logic_vector(17 downto 0); 
    of_x0: out std_logic
  );
end conv1_entity_11637058ac;

architecture structural of conv1_entity_11637058ac is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal all_0s_y_net: std_logic;
  signal all_1s_y_net: std_logic;
  signal and_y_net_x0: std_logic;
  signal ce_1_sg_x61: std_logic;
  signal clk_1_sg_x61: std_logic;
  signal invert1_op_net: std_logic;
  signal invert2_op_net: std_logic;
  signal invert3_op_net: std_logic;
  signal reinterpret4_output_port_net_x1: std_logic_vector(20 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic;
  signal slice3_y_net: std_logic;

begin
  ce_1_sg_x61 <= ce_1;
  clk_1_sg_x61 <= clk_1;
  reinterpret4_output_port_net_x1 <= din;
  dout <= adder_s_net_x5;
  of_x0 <= and_y_net_x0;

  all_0s: entity work.logical_3013ab8805
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      d0(0) => invert1_op_net,
      d1(0) => invert2_op_net,
      d2(0) => invert3_op_net,
      y(0) => all_0s_y_net
    );

  all_1s: entity work.logical_3013ab8805
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      d0(0) => slice1_y_net,
      d1(0) => slice2_y_net,
      d2(0) => slice3_y_net,
      y(0) => all_1s_y_net
    );

  and_x0: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => all_0s_y_net,
      d1(0) => all_1s_y_net,
      y(0) => and_y_net_x0
    );

  convert_f7847c8c42: entity work.convert_entity_f7847c8c42
    port map (
      ce_1 => ce_1_sg_x61,
      clk_1 => clk_1_sg_x61,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  invert1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      ip(0) => slice1_y_net,
      op(0) => invert1_op_net
    );

  invert2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      ip(0) => slice2_y_net,
      op(0) => invert2_op_net
    );

  invert3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      ip(0) => slice3_y_net,
      op(0) => invert3_op_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 20,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 19,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 18,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice3_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_convert/debus"

entity debus_entity_5fd018da5c is
  port (
    bus_in: in std_logic_vector(83 downto 0); 
    lsb_out1: out std_logic_vector(20 downto 0); 
    msb_out4: out std_logic_vector(20 downto 0); 
    out2: out std_logic_vector(20 downto 0); 
    out3: out std_logic_vector(20 downto 0)
  );
end debus_entity_5fd018da5c;

architecture structural of debus_entity_5fd018da5c is
  signal mux_y_net_x0: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(20 downto 0);
  signal slice1_y_net: std_logic_vector(20 downto 0);
  signal slice2_y_net: std_logic_vector(20 downto 0);
  signal slice3_y_net: std_logic_vector(20 downto 0);
  signal slice4_y_net: std_logic_vector(20 downto 0);

begin
  mux_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out4 <= reinterpret4_output_port_net_x2;
  out2 <= reinterpret2_output_port_net_x2;
  out3 <= reinterpret3_output_port_net_x2;

  reinterpret1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  reinterpret3: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x2
    );

  reinterpret4: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 20,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => mux_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 21,
      new_msb => 41,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => mux_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 42,
      new_msb => 62,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => mux_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 63,
      new_msb => 83,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => mux_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_convert"

entity bus_convert_entity_b21c3d5983 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(83 downto 0); 
    dout: out std_logic_vector(71 downto 0); 
    overflow: out std_logic_vector(3 downto 0)
  );
end bus_convert_entity_b21c3d5983;

architecture structural of bus_convert_entity_b21c3d5983 is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal adder_s_net_x8: std_logic_vector(17 downto 0);
  signal and_y_net_x4: std_logic;
  signal and_y_net_x5: std_logic;
  signal and_y_net_x6: std_logic;
  signal and_y_net_x7: std_logic;
  signal ce_1_sg_x68: std_logic;
  signal clk_1_sg_x68: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(3 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(20 downto 0);

begin
  ce_1_sg_x68 <= ce_1;
  clk_1_sg_x68 <= clk_1;
  mux_y_net_x1 <= din;
  dout <= concatenate_y_net_x2;
  overflow <= concatenate_y_net_x3;

  bussify_81a3739e19: entity work.bussify_entity_1d06622102
    port map (
      in1 => adder_s_net_x5,
      in2 => adder_s_net_x6,
      in3 => adder_s_net_x7,
      in4 => adder_s_net_x8,
      bus_out => concatenate_y_net_x2
    );

  conv1_11637058ac: entity work.conv1_entity_11637058ac
    port map (
      ce_1 => ce_1_sg_x68,
      clk_1 => clk_1_sg_x68,
      din => reinterpret4_output_port_net_x2,
      dout => adder_s_net_x5,
      of_x0 => and_y_net_x4
    );

  conv2_783611094b: entity work.conv1_entity_11637058ac
    port map (
      ce_1 => ce_1_sg_x68,
      clk_1 => clk_1_sg_x68,
      din => reinterpret3_output_port_net_x2,
      dout => adder_s_net_x6,
      of_x0 => and_y_net_x5
    );

  conv3_e0e7d86625: entity work.conv1_entity_11637058ac
    port map (
      ce_1 => ce_1_sg_x68,
      clk_1 => clk_1_sg_x68,
      din => reinterpret2_output_port_net_x2,
      dout => adder_s_net_x7,
      of_x0 => and_y_net_x6
    );

  conv4_4e5f30fb95: entity work.conv1_entity_11637058ac
    port map (
      ce_1 => ce_1_sg_x68,
      clk_1 => clk_1_sg_x68,
      din => reinterpret1_output_port_net_x2,
      dout => adder_s_net_x8,
      of_x0 => and_y_net_x7
    );

  debus_5fd018da5c: entity work.debus_entity_5fd018da5c
    port map (
      bus_in => mux_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

  of_bussify_c0a9d2e3fd: entity work.of_bussify_entity_be16087e66
    port map (
      in1 => and_y_net_x4,
      in2 => and_y_net_x5,
      in3 => and_y_net_x6,
      in4 => and_y_net_x7,
      bus_out => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_norm0/bussify"

entity bussify_entity_aa55880c0f is
  port (
    in1: in std_logic_vector(20 downto 0); 
    in2: in std_logic_vector(20 downto 0); 
    in3: in std_logic_vector(20 downto 0); 
    in4: in std_logic_vector(20 downto 0); 
    bus_out: out std_logic_vector(83 downto 0)
  );
end bussify_entity_aa55880c0f;

architecture structural of bussify_entity_aa55880c0f is
  signal concatenate_y_net_x0: std_logic_vector(83 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(20 downto 0);

begin
  conv1_dout_net_x0 <= in1;
  conv2_dout_net_x0 <= in2;
  conv3_dout_net_x0 <= in3;
  conv4_dout_net_x0 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_356a264444
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv1_dout_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv2_dout_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv3_dout_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv4_dout_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_norm0/debus"

entity debus_entity_3b6fb3cfa9 is
  port (
    bus_in: in std_logic_vector(79 downto 0); 
    lsb_out1: out std_logic_vector(19 downto 0); 
    msb_out4: out std_logic_vector(19 downto 0); 
    out2: out std_logic_vector(19 downto 0); 
    out3: out std_logic_vector(19 downto 0)
  );
end debus_entity_3b6fb3cfa9;

architecture structural of debus_entity_3b6fb3cfa9 is
  signal concat_y_net_x0: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic_vector(19 downto 0);
  signal slice2_y_net: std_logic_vector(19 downto 0);
  signal slice3_y_net: std_logic_vector(19 downto 0);
  signal slice4_y_net: std_logic_vector(19 downto 0);

begin
  concat_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 19,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 39,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 59,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 79,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_norm0"

entity bus_norm0_entity_19ac017aaf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(83 downto 0)
  );
end bus_norm0_entity_19ac017aaf;

architecture structural of bus_norm0_entity_19ac017aaf is
  signal ce_1_sg_x69: std_logic;
  signal clk_1_sg_x69: std_logic;
  signal concat_y_net_x1: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x69 <= ce_1;
  clk_1_sg_x69 <= clk_1;
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x1;

  bussify_aa55880c0f: entity work.bussify_entity_aa55880c0f
    port map (
      in1 => conv1_dout_net_x0,
      in2 => conv2_dout_net_x0,
      in3 => conv3_dout_net_x0,
      in4 => conv4_dout_net_x0,
      bus_out => concatenate_y_net_x1
    );

  conv1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x69,
      clk => clk_1_sg_x69,
      clr => '0',
      din => reinterpret4_output_port_net_x0,
      en => "1",
      dout => conv1_dout_net_x0
    );

  conv2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x69,
      clk => clk_1_sg_x69,
      clr => '0',
      din => reinterpret3_output_port_net_x0,
      en => "1",
      dout => conv2_dout_net_x0
    );

  conv3: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x69,
      clk => clk_1_sg_x69,
      clr => '0',
      din => reinterpret2_output_port_net_x0,
      en => "1",
      dout => conv3_dout_net_x0
    );

  conv4: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x69,
      clk => clk_1_sg_x69,
      clr => '0',
      din => reinterpret1_output_port_net_x0,
      en => "1",
      dout => conv4_dout_net_x0
    );

  debus_3b6fb3cfa9: entity work.debus_entity_3b6fb3cfa9
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_norm1/conv1"

entity conv1_entity_cfee4ad61e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(19 downto 0); 
    out_x0: out std_logic_vector(20 downto 0)
  );
end conv1_entity_cfee4ad61e;

architecture structural of conv1_entity_cfee4ad61e is
  signal adder_s_net_x4: std_logic_vector(20 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x70: std_logic;
  signal clk_1_sg_x70: std_logic;
  signal concat_y_net: std_logic_vector(20 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(20 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(19 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x70 <= ce_1;
  clk_1_sg_x70 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.addsub_43b12feb7d
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x70,
      clk => clk_1_sg_x70,
      clr => '0',
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_b366689086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_c615d93998
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_b1e9d7c303
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_norm1"

entity bus_norm1_entity_d801aceba7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(83 downto 0)
  );
end bus_norm1_entity_d801aceba7;

architecture structural of bus_norm1_entity_d801aceba7 is
  signal adder_s_net_x4: std_logic_vector(20 downto 0);
  signal adder_s_net_x5: std_logic_vector(20 downto 0);
  signal adder_s_net_x6: std_logic_vector(20 downto 0);
  signal adder_s_net_x7: std_logic_vector(20 downto 0);
  signal ce_1_sg_x74: std_logic;
  signal clk_1_sg_x74: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x74 <= ce_1;
  clk_1_sg_x74 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_c819990780: entity work.bussify_entity_aa55880c0f
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_cfee4ad61e: entity work.conv1_entity_cfee4ad61e
    port map (
      ce_1 => ce_1_sg_x74,
      clk_1 => clk_1_sg_x74,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_aaf233eaa8: entity work.conv1_entity_cfee4ad61e
    port map (
      ce_1 => ce_1_sg_x74,
      clk_1 => clk_1_sg_x74,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_4b74605deb: entity work.conv1_entity_cfee4ad61e
    port map (
      ce_1 => ce_1_sg_x74,
      clk_1 => clk_1_sg_x74,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_4111a03a03: entity work.conv1_entity_cfee4ad61e
    port map (
      ce_1 => ce_1_sg_x74,
      clk_1 => clk_1_sg_x74,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_fdd218b3f9: entity work.debus_entity_71deb38b98
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_scale"

entity bus_scale_entity_cc780061b4 is
  port (
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_scale_entity_cc780061b4;

architecture structural of bus_scale_entity_cc780061b4 is
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal scale1_op_net_x0: std_logic_vector(19 downto 0);
  signal scale2_op_net_x0: std_logic_vector(19 downto 0);
  signal scale3_op_net_x0: std_logic_vector(19 downto 0);
  signal scale4_op_net_x0: std_logic_vector(19 downto 0);

begin
  concat_y_net_x3 <= din;
  dout <= concatenate_y_net_x4;

  bussify_76471ddda6: entity work.bussify_entity_6546069b97
    port map (
      in1 => scale1_op_net_x0,
      in2 => scale2_op_net_x0,
      in3 => scale3_op_net_x0,
      in4 => scale4_op_net_x0,
      bus_out => concatenate_y_net_x4
    );

  debus_37f472a9a7: entity work.debus_entity_3b6fb3cfa9
    port map (
      bus_in => concat_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  scale1: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret4_output_port_net_x0,
      op => scale1_op_net_x0
    );

  scale2: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret3_output_port_net_x0,
      op => scale2_op_net_x0
    );

  scale3: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret2_output_port_net_x0,
      op => scale3_op_net_x0
    );

  scale4: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret1_output_port_net_x0,
      op => scale4_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/bus_sub"

entity bus_sub_entity_5f1ccce5f7 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(37 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(39 downto 0)
  );
end bus_sub_entity_5f1ccce5f7;

architecture structural of bus_sub_entity_5f1ccce5f7 is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal ce_1_sg_x75: std_logic;
  signal clk_1_sg_x75: std_logic;
  signal concatenate_y_net_x4: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  reinterpret1_output_port_net_x5 <= a;
  concatenate_y_net_x4 <= b;
  ce_1_sg_x75 <= ce_1;
  clk_1_sg_x75 <= clk_1;
  dout <= concatenate_y_net_x5;

  a_debus_6b1eb6941c: entity work.a_debus_entity_c0242f8ce0
    port map (
      bus_in => reinterpret1_output_port_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_a0497faccc62b6b2",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x75,
      clk => clk_1_sg_x75,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_a0497faccc62b6b2",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x75,
      clk => clk_1_sg_x75,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_52927e5641: entity work.b_debus_entity_98717e8269
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_b2e31fcc70: entity work.op_bussify_entity_f21ce432ef
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert/conv1"

entity conv1_entity_88c6c6d96e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(36 downto 0); 
    out_x0: out std_logic_vector(18 downto 0)
  );
end conv1_entity_88c6c6d96e;

architecture structural of conv1_entity_88c6c6d96e is
  signal adder_s_net_x2: std_logic_vector(18 downto 0);
  signal almost_half_op_net: std_logic_vector(34 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x76: std_logic;
  signal clk_1_sg_x76: std_logic;
  signal concat_y_net: std_logic_vector(37 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(37 downto 0);
  signal force2_output_port_net: std_logic_vector(34 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(36 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(36 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x76 <= ce_1;
  clk_1_sg_x76 <= clk_1;
  reinterpret2_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x2;

  adder: entity work.addsub_82254b26db
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      s => adder_s_net_x2
    );

  almost_half: entity work.constant_2da6af93c2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 36,
      x_width => 37,
      y_width => 1
    )
    port map (
      x => reinterpret2_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_83820b2faf
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_620dd01637
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_ec14c62a89
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert/debus"

entity debus_entity_f1c09f94b9 is
  port (
    bus_in: in std_logic_vector(73 downto 0); 
    lsb_out1: out std_logic_vector(36 downto 0); 
    msb_out2: out std_logic_vector(36 downto 0)
  );
end debus_entity_f1c09f94b9;

architecture structural of debus_entity_f1c09f94b9 is
  signal reinterpret1_output_port_net_x1: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(36 downto 0);
  signal slice1_y_net: std_logic_vector(36 downto 0);
  signal slice2_y_net: std_logic_vector(36 downto 0);

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out2 <= reinterpret2_output_port_net_x1;

  reinterpret1: entity work.reinterpret_5b4829fb41
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_5b4829fb41
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 36,
      x_width => 74,
      y_width => 37
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 37,
      new_msb => 73,
      x_width => 74,
      y_width => 37
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert"

entity bus_convert_entity_a82e0e1650 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(73 downto 0); 
    misci: in std_logic_vector(36 downto 0); 
    dout: out std_logic_vector(37 downto 0); 
    misco: out std_logic_vector(36 downto 0)
  );
end bus_convert_entity_a82e0e1650;

architecture structural of bus_convert_entity_a82e0e1650 is
  signal adder_s_net_x2: std_logic_vector(18 downto 0);
  signal adder_s_net_x3: std_logic_vector(18 downto 0);
  signal ce_1_sg_x78: std_logic;
  signal clk_1_sg_x78: std_logic;
  signal concatenate_y_net_x6: std_logic_vector(37 downto 0);
  signal dmisc_q_net_x1: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(36 downto 0);

begin
  ce_1_sg_x78 <= ce_1;
  clk_1_sg_x78 <= clk_1;
  reinterpret1_output_port_net_x3 <= din;
  dmisc_q_net_x1 <= misci;
  dout <= concatenate_y_net_x6;
  misco <= dmisc_q_net_x2;

  bussify_91f9dbc7f3: entity work.op_bussify_entity_8ee3422350
    port map (
      in1 => adder_s_net_x2,
      in2 => adder_s_net_x3,
      bus_out => concatenate_y_net_x6
    );

  conv1_88c6c6d96e: entity work.conv1_entity_88c6c6d96e
    port map (
      ce_1 => ce_1_sg_x78,
      clk_1 => clk_1_sg_x78,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x2
    );

  conv2_937900189b: entity work.conv1_entity_88c6c6d96e
    port map (
      ce_1 => ce_1_sg_x78,
      clk_1 => clk_1_sg_x78,
      in_x0 => reinterpret1_output_port_net_x2,
      out_x0 => adder_s_net_x3
    );

  debus_f1c09f94b9: entity work.debus_entity_f1c09f94b9
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  dmisc: entity work.delay_64530ed2c8
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      d => dmisc_q_net_x1,
      q => dmisc_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_create"

entity bus_create_entity_9c2c0dccf0 is
  port (
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic; 
    in3: in std_logic_vector(35 downto 0); 
    bus_out: out std_logic_vector(72 downto 0)
  );
end bus_create_entity_9c2c0dccf0;

architecture structural of bus_create_entity_9c2c0dccf0 is
  signal concatenate_y_net_x0: std_logic_vector(72 downto 0);
  signal delay_q_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic_vector(35 downto 0);

begin
  mux_y_net_x1 <= in1;
  mux_y_net_x2 <= in2;
  delay_q_net_x0 <= in3;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_b28df1ab2e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x1,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => mux_y_net_x2,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => delay_q_net_x0,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_expand"

entity bus_expand_entity_ad772b3d60 is
  port (
    bus_in: in std_logic_vector(72 downto 0); 
    lsb_out1: out std_logic_vector(36 downto 0); 
    msb_out2: out std_logic_vector(35 downto 0)
  );
end bus_expand_entity_ad772b3d60;

architecture structural of bus_expand_entity_ad772b3d60 is
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(36 downto 0);
  signal slice2_y_net: std_logic_vector(35 downto 0);

begin
  delay1_q_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_892b735f0d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 36,
      x_width => 73,
      y_width => 37
    )
    port map (
      x => delay1_q_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 37,
      new_msb => 72,
      x_width => 73,
      y_width => 36
    )
    port map (
      x => delay1_q_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_expand1"

entity bus_expand1_entity_e394667c48 is
  port (
    bus_in: in std_logic_vector(36 downto 0); 
    lsb_out1: out std_logic_vector(35 downto 0); 
    msb_out2: out std_logic
  );
end bus_expand1_entity_e394667c48;

architecture structural of bus_expand1_entity_e394667c48 is
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);
  signal slice2_y_net_x0: std_logic;

begin
  dmisc_q_net_x3 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x6;
  msb_out2 <= slice2_y_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x6
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 37,
      y_width => 36
    )
    port map (
      x => dmisc_q_net_x3,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 36,
      x_width => 37,
      y_width => 1
    )
    port map (
      x => dmisc_q_net_x3,
      y(0) => slice2_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/a*b_bussify"

entity a_b_bussify_entity_2a7d6fa717 is
  port (
    in1: in std_logic_vector(73 downto 0); 
    bus_out: out std_logic_vector(73 downto 0)
  );
end a_b_bussify_entity_2a7d6fa717;

architecture structural of a_b_bussify_entity_2a7d6fa717 is
  signal concat_y_net_x0: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(73 downto 0);

begin
  concat_y_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x4;

  reinterpret1: entity work.reinterpret_efdf1c3890
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net_x0,
      output_port => reinterpret1_output_port_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/a_debus"

entity a_debus_entity_9378c272e1 is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    msb_lsb_out1: out std_logic_vector(35 downto 0)
  );
end a_debus_entity_9378c272e1;

architecture structural of a_debus_entity_9378c272e1 is
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 36,
      y_width => 36
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/c_to_ri"

entity c_to_ri_entity_8f95d0368d is
  port (
    c: in std_logic_vector(35 downto 0); 
    im: out std_logic_vector(17 downto 0); 
    re: out std_logic_vector(17 downto 0)
  );
end c_to_ri_entity_8f95d0368d;

architecture structural of c_to_ri_entity_8f95d0368d is
  signal force_im_output_port_net_x0: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice_im_y_net: std_logic_vector(17 downto 0);
  signal slice_re_y_net: std_logic_vector(17 downto 0);

begin
  reinterpret1_output_port_net_x3 <= c;
  im <= force_im_output_port_net_x0;
  re <= force_re_output_port_net_x0;

  force_im: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_im_y_net,
      output_port => force_im_output_port_net_x0
    );

  force_re: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_re_y_net,
      output_port => force_re_output_port_net_x0
    );

  slice_im: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret1_output_port_net_x3,
      y => slice_im_y_net
    );

  slice_re: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret1_output_port_net_x3,
      y => slice_re_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/ri_to_c"

entity ri_to_c_entity_8792409687 is
  port (
    im: in std_logic_vector(36 downto 0); 
    re: in std_logic_vector(36 downto 0); 
    c: out std_logic_vector(73 downto 0)
  );
end ri_to_c_entity_8792409687;

architecture structural of ri_to_c_entity_8792409687 is
  signal concat_y_net_x1: std_logic_vector(73 downto 0);
  signal convert_im_dout_net_x0: std_logic_vector(36 downto 0);
  signal convert_re_dout_net_x0: std_logic_vector(36 downto 0);
  signal force_im_output_port_net: std_logic_vector(36 downto 0);
  signal force_re_output_port_net: std_logic_vector(36 downto 0);

begin
  convert_im_dout_net_x0 <= im;
  convert_re_dout_net_x0 <= re;
  c <= concat_y_net_x1;

  concat: entity work.concat_56d57d2c92
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x1
    );

  force_im: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_im_dout_net_x0,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_re_dout_net_x0,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1"

entity mult1_entity_c9146ccfd6 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ab: out std_logic_vector(73 downto 0)
  );
end mult1_entity_c9146ccfd6;

architecture structural of mult1_entity_c9146ccfd6 is
  signal addsub_im_s_net: std_logic_vector(36 downto 0);
  signal addsub_re_s_net: std_logic_vector(36 downto 0);
  signal ce_1_sg_x79: std_logic;
  signal clk_1_sg_x79: std_logic;
  signal concat_y_net_x2: std_logic_vector(73 downto 0);
  signal convert_im_dout_net_x0: std_logic_vector(36 downto 0);
  signal convert_re_dout_net_x0: std_logic_vector(36 downto 0);
  signal force_im_output_port_net_x0: std_logic_vector(17 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x0: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal imim_p_net: std_logic_vector(35 downto 0);
  signal imre_p_net: std_logic_vector(35 downto 0);
  signal reim_p_net: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal rere_p_net: std_logic_vector(35 downto 0);

begin
  reinterpret1_output_port_net_x5 <= a;
  reinterpret1_output_port_net_x6 <= b;
  ce_1_sg_x79 <= ce_1;
  clk_1_sg_x79 <= clk_1;
  ab <= concat_y_net_x2;

  addsub_im: entity work.addsub_4ded11ba54
    port map (
      a => imre_p_net,
      b => reim_p_net,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      s => addsub_im_s_net
    );

  addsub_re: entity work.addsub_8dd4a43ef5
    port map (
      a => rere_p_net,
      b => imim_p_net,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      s => addsub_re_s_net
    );

  c_to_ri1_6f24614ac7: entity work.c_to_ri_entity_8f95d0368d
    port map (
      c => reinterpret1_output_port_net_x6,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  c_to_ri_8f95d0368d: entity work.c_to_ri_entity_8f95d0368d
    port map (
      c => reinterpret1_output_port_net_x5,
      im => force_im_output_port_net_x0,
      re => force_re_output_port_net_x0
    );

  convert_im: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 34,
      din_width => 37,
      dout_arith => 2,
      dout_bin_pt => 34,
      dout_width => 37,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      din => addsub_im_s_net,
      en => "1",
      dout => convert_im_dout_net_x0
    );

  convert_re: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 34,
      din_width => 37,
      dout_arith => 2,
      dout_bin_pt => 34,
      dout_width => 37,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      din => addsub_re_s_net,
      en => "1",
      dout => convert_re_dout_net_x0
    );

  imim: entity work.mult_f295e5f0f2
    port map (
      a => force_im_output_port_net_x0,
      b => force_im_output_port_net_x1,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      p => imim_p_net
    );

  imre: entity work.mult_f295e5f0f2
    port map (
      a => force_im_output_port_net_x0,
      b => force_re_output_port_net_x1,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      p => imre_p_net
    );

  reim: entity work.mult_f295e5f0f2
    port map (
      a => force_re_output_port_net_x0,
      b => force_im_output_port_net_x1,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      p => reim_p_net
    );

  rere: entity work.mult_f295e5f0f2
    port map (
      a => force_re_output_port_net_x0,
      b => force_re_output_port_net_x1,
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      clr => '0',
      p => rere_p_net
    );

  ri_to_c_8792409687: entity work.ri_to_c_entity_8792409687
    port map (
      im => convert_im_dout_net_x0,
      re => convert_re_dout_net_x0,
      c => concat_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/repa/bussify"

entity bussify_entity_d6ea8ebb9b is
  port (
    in1: in std_logic_vector(35 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end bussify_entity_d6ea8ebb9b;

architecture structural of bussify_entity_d6ea8ebb9b is
  signal register0_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  register0_q_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => register0_q_net_x0,
      output_port => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/repa/din1"

entity din1_entity_080142ebc1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic_vector(35 downto 0); 
    q: out std_logic_vector(35 downto 0)
  );
end din1_entity_080142ebc1;

architecture structural of din1_entity_080142ebc1 is
  signal ce_1_sg_x80: std_logic;
  signal clk_1_sg_x80: std_logic;
  signal concat_y_net_x0: std_logic_vector(35 downto 0);
  signal register0_q_net_x1: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x80 <= ce_1;
  clk_1_sg_x80 <= clk_1;
  concat_y_net_x0 <= d;
  q <= register0_q_net_x1;

  register0: entity work.xlregister
    generic map (
      d_width => 36,
      init_value => b"000000000000000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x80,
      clk => clk_1_sg_x80,
      d => concat_y_net_x0,
      en => "1",
      rst => "0",
      q => register0_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/repa"

entity repa_entity_9388816dba is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(35 downto 0); 
    out_x0: out std_logic_vector(35 downto 0)
  );
end repa_entity_9388816dba;

architecture structural of repa_entity_9388816dba is
  signal ce_1_sg_x81: std_logic;
  signal clk_1_sg_x81: std_logic;
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal register0_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x81 <= ce_1;
  clk_1_sg_x81 <= clk_1;
  concat_y_net_x1 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x3;

  bussify_d6ea8ebb9b: entity work.bussify_entity_d6ea8ebb9b
    port map (
      in1 => register0_q_net_x1,
      bus_out => reinterpret1_output_port_net_x3
    );

  din1_080142ebc1: entity work.din1_entity_080142ebc1
    port map (
      ce_1 => ce_1_sg_x81,
      clk_1 => clk_1_sg_x81,
      d => concat_y_net_x1,
      q => register0_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult"

entity bus_mult_entity_f9d9d4b2f7 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(36 downto 0); 
    a_b: out std_logic_vector(73 downto 0); 
    misco: out std_logic_vector(36 downto 0)
  );
end bus_mult_entity_f9d9d4b2f7;

architecture structural of bus_mult_entity_f9d9d4b2f7 is
  signal ce_1_sg_x84: std_logic;
  signal clk_1_sg_x84: std_logic;
  signal concat_y_net_x2: std_logic_vector(73 downto 0);
  signal concat_y_net_x3: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);

begin
  concat_y_net_x3 <= a;
  reinterpret2_output_port_net_x3 <= b;
  ce_1_sg_x84 <= ce_1;
  clk_1_sg_x84 <= clk_1;
  reinterpret1_output_port_net_x8 <= misci;
  a_b <= reinterpret1_output_port_net_x9;
  misco <= dmisc_q_net_x2;

  a_b_bussify_2a7d6fa717: entity work.a_b_bussify_entity_2a7d6fa717
    port map (
      in1 => concat_y_net_x2,
      bus_out => reinterpret1_output_port_net_x9
    );

  a_debus_9378c272e1: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x5
    );

  b_debus_64000166bd: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => reinterpret1_output_port_net_x7,
      msb_lsb_out1 => reinterpret1_output_port_net_x6
    );

  dmisc: entity work.delay_2d0f74b2c1
    port map (
      ce => ce_1_sg_x84,
      clk => clk_1_sg_x84,
      clr => '0',
      d => reinterpret1_output_port_net_x8,
      q => dmisc_q_net_x2
    );

  mult1_c9146ccfd6: entity work.mult1_entity_c9146ccfd6
    port map (
      a => reinterpret1_output_port_net_x5,
      b => reinterpret1_output_port_net_x6,
      ce_1 => ce_1_sg_x84,
      clk_1 => clk_1_sg_x84,
      ab => concat_y_net_x2
    );

  repa_9388816dba: entity work.repa_entity_9388816dba
    port map (
      ce_1 => ce_1_sg_x84,
      clk_1 => clk_1_sg_x84,
      in_x0 => concat_y_net_x3,
      out_x0 => reinterpret1_output_port_net_x3
    );

  repb_41919bcfb1: entity work.repa_entity_9388816dba
    port map (
      ce_1 => ce_1_sg_x84,
      clk_1 => clk_1_sg_x84,
      in_x0 => reinterpret2_output_port_net_x3,
      out_x0 => reinterpret1_output_port_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_2af7d3a329 is
  port (
    in_x0: in std_logic_vector(8 downto 0); 
    out_x0: out std_logic_vector(8 downto 0)
  );
end bit_reverse_entity_2af7d3a329;

architecture structural of bit_reverse_entity_2af7d3a329 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(8 downto 0);
  signal slice_y_net_x0: std_logic_vector(8 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  concat: entity work.concat_0cc72cd991
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_b94e068100 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(8 downto 0); 
    add: out std_logic_vector(8 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_b94e068100;

architecture structural of add_convert0_entity_b94e068100 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(8 downto 0);
  signal ce_1_sg_x85: std_logic;
  signal clk_1_sg_x85: std_logic;
  signal concat_y_net: std_logic_vector(9 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal delay13_q_net: std_logic_vector(8 downto 0);
  signal delay14_q_net: std_logic_vector(8 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(9 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(7 downto 0);
  signal new_add_y_net: std_logic_vector(8 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x85 <= ce_1;
  clk_1_sg_x85 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_7eef56098d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 9,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 9,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_09771002d6
    port map (
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_09771002d6
    port map (
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x85,
      clk => clk_1_sg_x85,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9779a5cf83
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 10,
      y_width => 8
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 10,
      y_width => 9
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 9,
      x_width => 10,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_743220f083 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(8 downto 0); 
    add: out std_logic_vector(8 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_743220f083;

architecture structural of add_convert1_entity_743220f083 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x86: std_logic;
  signal clk_1_sg_x86: std_logic;
  signal concat_y_net: std_logic_vector(9 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal delay13_q_net: std_logic_vector(8 downto 0);
  signal delay14_q_net: std_logic_vector(8 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(9 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(7 downto 0);
  signal new_add_y_net: std_logic_vector(8 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x86 <= ce_1;
  clk_1_sg_x86 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_7eef56098d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 9,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 9,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_09771002d6
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_09771002d6
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9779a5cf83
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 10,
      y_width => 8
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 10,
      y_width => 9
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 9,
      x_width => 10,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/invert0"

entity invert0_entity_e94ce56a25 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(17 downto 0); 
    negate_x0: in std_logic; 
    out_x0: out std_logic_vector(17 downto 0)
  );
end invert0_entity_e94ce56a25;

architecture structural of invert0_entity_e94ce56a25 is
  signal ce_1_sg_x87: std_logic;
  signal clk_1_sg_x87: std_logic;
  signal delay10_q_net_x0: std_logic;
  signal delay20_q_net: std_logic_vector(17 downto 0);
  signal delay21_q_net: std_logic;
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x0: std_logic_vector(17 downto 0);
  signal negate_op_net: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x87 <= ce_1;
  clk_1_sg_x87 <= clk_1;
  lookup_douta_net_x0 <= in_x0;
  delay10_q_net_x0 <= negate_x0;
  out_x0 <= mux_y_net_x0;

  delay20: entity work.delay_b6092ad150
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      d => lookup_douta_net_x0,
      q => delay20_q_net
    );

  delay21: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      d(0) => delay10_q_net_x0,
      q(0) => delay21_q_net
    );

  mux: entity work.mux_bc64561e19
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      d0 => delay20_q_net,
      d1 => negate_op_net,
      sel(0) => delay21_q_net,
      y => mux_y_net_x0
    );

  negate: entity work.negate_206b7f76d8
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      ip => lookup_douta_net_x0,
      op => negate_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/invert1"

entity invert1_entity_56100eb48e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(17 downto 0); 
    misci: in std_logic_vector(72 downto 0); 
    negate_x0: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end invert1_entity_56100eb48e;

architecture structural of invert1_entity_56100eb48e is
  signal ce_1_sg_x88: std_logic;
  signal clk_1_sg_x88: std_logic;
  signal delay1_q_net_x1: std_logic_vector(72 downto 0);
  signal delay20_q_net: std_logic_vector(17 downto 0);
  signal delay21_q_net: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x0: std_logic_vector(17 downto 0);
  signal negate_op_net: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x88 <= ce_1;
  clk_1_sg_x88 <= clk_1;
  lookup_doutb_net_x0 <= in_x0;
  delay_q_net_x0 <= misci;
  delay8_q_net_x0 <= negate_x0;
  misco <= delay1_q_net_x1;
  out_x0 <= mux_y_net_x0;

  delay1: entity work.delay_7097453b2c
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d => delay_q_net_x0,
      q => delay1_q_net_x1
    );

  delay20: entity work.delay_b6092ad150
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d => lookup_doutb_net_x0,
      q => delay20_q_net
    );

  delay21: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d(0) => delay8_q_net_x0,
      q(0) => delay21_q_net
    );

  mux: entity work.mux_bc64561e19
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d0 => delay20_q_net,
      d1 => negate_op_net,
      sel(0) => delay21_q_net,
      y => mux_y_net_x0
    );

  negate: entity work.negate_206b7f76d8
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      ip => lookup_doutb_net_x0,
      op => negate_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_4c5f50bca4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(8 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_4c5f50bca4;

architecture structural of cosin_entity_4c5f50bca4 is
  signal assert_dout_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x89: std_logic;
  signal clk_1_sg_x89: std_logic;
  signal concat_y_net_x1: std_logic_vector(8 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(8 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x89 <= ce_1;
  clk_1_sg_x89 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_b94e068100: entity work.add_convert0_entity_b94e068100
    port map (
      ce_1 => ce_1_sg_x89,
      clk_1 => clk_1_sg_x89,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_743220f083: entity work.add_convert1_entity_743220f083
    port map (
      ce_1 => ce_1_sg_x89,
      clk_1 => clk_1_sg_x89,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 9,
      dout_width => 9
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x89,
      clk => clk_1_sg_x89,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x89,
      clk => clk_1_sg_x89,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x89,
      clk => clk_1_sg_x89,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_e94ce56a25: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x89,
      clk_1 => clk_1_sg_x89,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_56100eb48e: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x89,
      clk_1 => clk_1_sg_x89,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_core
    generic map (
      c_address_width_a => 9,
      c_address_width_b => 9,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_c1a8b20e2e422729",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x89,
      a_clk => clk_1_sg_x89,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x89,
      b_clk => clk_1_sg_x89,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/ri_to_c"

entity ri_to_c_entity_7d26fbf4c5 is
  port (
    im: in std_logic_vector(17 downto 0); 
    re: in std_logic_vector(17 downto 0); 
    c: out std_logic_vector(35 downto 0)
  );
end ri_to_c_entity_7d26fbf4c5;

architecture structural of ri_to_c_entity_7d26fbf4c5 is
  signal concat_y_net_x4: std_logic_vector(35 downto 0);
  signal force_im_output_port_net: std_logic_vector(17 downto 0);
  signal force_re_output_port_net: std_logic_vector(17 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);

begin
  mux_y_net_x5 <= im;
  mux_y_net_x4 <= re;
  c <= concat_y_net_x4;

  concat: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x4
    );

  force_im: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x5,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x4,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_0c3bb01e4d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_0c3bb01e4d;

architecture structural of coeff_gen_entity_0c3bb01e4d is
  signal ce_1_sg_x90: std_logic;
  signal clk_1_sg_x90: std_logic;
  signal concat_y_net_x1: std_logic_vector(8 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(8 downto 0);

begin
  ce_1_sg_x90 <= ce_1;
  clk_1_sg_x90 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_2af7d3a329: entity work.bit_reverse_entity_2af7d3a329
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_4c5f50bca4: entity work.cosin_entity_4c5f50bca4
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_7d26fbf4c5: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 11,
      x_width => 12,
      y_width => 9
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct/twiddle"

entity twiddle_entity_d1767287eb is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_d1767287eb;

architecture structural of twiddle_entity_d1767287eb is
  signal ce_1_sg_x91: std_logic;
  signal clk_1_sg_x91: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal delay_q_net_x1: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  delay_q_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x91 <= ce_1;
  clk_1_sg_x91 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_a82e0e1650: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x91,
      clk_1 => clk_1_sg_x91,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_9c2c0dccf0: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => delay_q_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_e394667c48: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_ad772b3d60: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_f9d9d4b2f7: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x91,
      clk_1 => clk_1_sg_x91,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_0c3bb01e4d: entity work.coeff_gen_entity_0c3bb01e4d
    port map (
      ce_1 => ce_1_sg_x91,
      clk_1 => clk_1_sg_x91,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/butterfly_direct"

entity butterfly_direct_entity_586c981496 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_586c981496;

architecture structural of butterfly_direct_entity_586c981496 is
  signal ce_1_sg_x92: std_logic;
  signal clk_1_sg_x92: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal delay_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  delay_q_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x92 <= ce_1;
  clk_1_sg_x92 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_fda2dbc1e4: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      dout => concatenate_y_net_x3
    );

  bus_convert_b21c3d5983: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_16b072c24d: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_19ac017aaf: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_d801aceba7: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_5d0abcce3e: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_cc780061b4: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_5f1ccce5f7: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x92,
      clk => clk_1_sg_x92,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x92,
      clk => clk_1_sg_x92,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_9c3e6d2a10: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x92,
      clk => clk_1_sg_x92,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_d1767287eb: entity work.twiddle_entity_d1767287eb
    port map (
      ai => delay_q_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x92,
      clk_1 => clk_1_sg_x92,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/delay_b"

entity delay_b_entity_bfead57ec1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_bfead57ec1;

architecture structural of delay_b_entity_bfead57ec1 is
  signal ce_1_sg_x93: std_logic;
  signal clk_1_sg_x93: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x93 <= ce_1;
  clk_1_sg_x93 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= delay_q_net_x3;

  delay: entity work.delay_faa52967c8
    port map (
      ce => ce_1_sg_x93,
      clk => clk_1_sg_x93,
      clr => '0',
      d => mux1_y_net_x0,
      q => delay_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10/sync_delay"

entity sync_delay_entity_93462c1816 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_93462c1816;

architecture structural of sync_delay_entity_93462c1816 is
  signal ce_1_sg_x95: std_logic;
  signal clk_1_sg_x95: std_logic;
  signal constant1_op_net: std_logic_vector(3 downto 0);
  signal constant2_op_net: std_logic_vector(3 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(3 downto 0);
  signal counter_op_net: std_logic_vector(3 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x95 <= ce_1;
  clk_1_sg_x95 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_145086465d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_67ad97ca70
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_a1505185555f1882",
      op_arith => xlUnsigned,
      op_width => 4
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_4d3cfceaf4
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_d930162434
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_10"

entity fft_stage_10_entity_3b39e0a900 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_10_entity_3b39e0a900;

architecture structural of fft_stage_10_entity_3b39e0a900 is
  signal ce_1_sg_x96: std_logic;
  signal clk_1_sg_x96: std_logic;
  signal counter_op_net: std_logic_vector(3 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal delay_q_net_x0: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal delay_q_net_x4: std_logic_vector(35 downto 0);
  signal fft_shift_net_x1: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x96 <= ce_1;
  clk_1_sg_x96 <= clk_1;
  reinterpret2_output_port_net_x0 <= in1;
  reinterpret1_output_port_net_x1 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x1 <= shift;
  delay0_q_net_x1 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x12;
  sync_out <= delay0_q_net_x2;

  butterfly_direct_586c981496: entity work.butterfly_direct_entity_586c981496
    port map (
      a => delay_q_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x96,
      clk_1 => clk_1_sg_x96,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x12,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x2
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_7789a80a5b2a8160",
      op_arith => xlUnsigned,
      op_width => 4
    )
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x1,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      d(0) => delay0_q_net_x1,
      q(0) => delay_q_net_x0
    );

  delay_b_bfead57ec1: entity work.delay_b_entity_bfead57ec1
    port map (
      ce_1 => ce_1_sg_x96,
      clk_1 => clk_1_sg_x96,
      din => mux1_y_net_x0,
      dout => delay_q_net_x3
    );

  delay_f_59a06da88c: entity work.delay_b_entity_bfead57ec1
    port map (
      ce_1 => ce_1_sg_x96,
      clk_1 => clk_1_sg_x96,
      din => reinterpret1_output_port_net_x1,
      dout => delay_q_net_x4
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      d0 => delay_q_net_x4,
      d1 => reinterpret2_output_port_net_x0,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      d0 => reinterpret2_output_port_net_x0,
      d1 => delay_q_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x1,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_93462c1816: entity work.sync_delay_entity_93462c1816
    port map (
      ce_1 => ce_1_sg_x96,
      clk_1 => clk_1_sg_x96,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_db36d4e0f5 is
  port (
    in_x0: in std_logic_vector(9 downto 0); 
    out_x0: out std_logic_vector(9 downto 0)
  );
end bit_reverse_entity_db36d4e0f5;

architecture structural of bit_reverse_entity_db36d4e0f5 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(9 downto 0);
  signal slice_y_net_x0: std_logic_vector(9 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_e774b32dc9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_db6a73eb6b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(9 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_db6a73eb6b;

architecture structural of add_convert0_entity_db6a73eb6b is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(9 downto 0);
  signal ce_1_sg_x123: std_logic;
  signal clk_1_sg_x123: std_logic;
  signal concat_y_net: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic_vector(9 downto 0);
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(10 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(8 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x123 <= ce_1;
  clk_1_sg_x123 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_4fd36a24a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 10,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_811dd91a3d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 11,
      y_width => 9
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 11,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 10,
      x_width => 11,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_1b4024ca70 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(9 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_1b4024ca70;

architecture structural of add_convert1_entity_1b4024ca70 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(9 downto 0);
  signal ce_1_sg_x124: std_logic;
  signal clk_1_sg_x124: std_logic;
  signal concat_y_net: std_logic_vector(10 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic_vector(9 downto 0);
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(10 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(8 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x124 <= ce_1;
  clk_1_sg_x124 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_4fd36a24a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 10,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x124,
      clk => clk_1_sg_x124,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_811dd91a3d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 11,
      y_width => 9
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 11,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 10,
      x_width => 11,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_65a50ac871 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(9 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_65a50ac871;

architecture structural of cosin_entity_65a50ac871 is
  signal assert_dout_net_x1: std_logic_vector(9 downto 0);
  signal ce_1_sg_x127: std_logic;
  signal clk_1_sg_x127: std_logic;
  signal concat_y_net_x1: std_logic_vector(9 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(9 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x127 <= ce_1;
  clk_1_sg_x127 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_db6a73eb6b: entity work.add_convert0_entity_db6a73eb6b
    port map (
      ce_1 => ce_1_sg_x127,
      clk_1 => clk_1_sg_x127,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_1b4024ca70: entity work.add_convert1_entity_1b4024ca70
    port map (
      ce_1 => ce_1_sg_x127,
      clk_1 => clk_1_sg_x127,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 10,
      dout_width => 10
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x127,
      clk => clk_1_sg_x127,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x127,
      clk => clk_1_sg_x127,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x127,
      clk => clk_1_sg_x127,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_f90c719cbc: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x127,
      clk_1 => clk_1_sg_x127,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_0cff7f13b2: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x127,
      clk_1 => clk_1_sg_x127,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_core
    generic map (
      c_address_width_a => 10,
      c_address_width_b => 10,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_9f585cf1e3329833",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x127,
      a_clk => clk_1_sg_x127,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x127,
      b_clk => clk_1_sg_x127,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_f755d375ac is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_f755d375ac;

architecture structural of coeff_gen_entity_f755d375ac is
  signal ce_1_sg_x128: std_logic;
  signal clk_1_sg_x128: std_logic;
  signal concat_y_net_x1: std_logic_vector(9 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x128 <= ce_1;
  clk_1_sg_x128 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_db36d4e0f5: entity work.bit_reverse_entity_db36d4e0f5
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_65a50ac871: entity work.cosin_entity_65a50ac871
    port map (
      ce_1 => ce_1_sg_x128,
      clk_1 => clk_1_sg_x128,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x128,
      clk => clk_1_sg_x128,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_7498c4690d: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 11,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct/twiddle"

entity twiddle_entity_e43eb2f177 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_e43eb2f177;

architecture structural of twiddle_entity_e43eb2f177 is
  signal ce_1_sg_x129: std_logic;
  signal clk_1_sg_x129: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal delay_q_net_x1: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  delay_q_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x129 <= ce_1;
  clk_1_sg_x129 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_e9bdbd1046: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x129,
      clk_1 => clk_1_sg_x129,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_6b84799eba: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => delay_q_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_64f8dfb179: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_d0b7647b56: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_c71dedf907: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x129,
      clk_1 => clk_1_sg_x129,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_f755d375ac: entity work.coeff_gen_entity_f755d375ac
    port map (
      ce_1 => ce_1_sg_x129,
      clk_1 => clk_1_sg_x129,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/butterfly_direct"

entity butterfly_direct_entity_6a735ce8e8 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_6a735ce8e8;

architecture structural of butterfly_direct_entity_6a735ce8e8 is
  signal ce_1_sg_x130: std_logic;
  signal clk_1_sg_x130: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal delay_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  delay_q_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x130 <= ce_1;
  clk_1_sg_x130 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_50d28544a9: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      dout => concatenate_y_net_x3
    );

  bus_convert_f7f638beba: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_3e3be77c79: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_706dadbee9: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_5fddbde300: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_4bcad4d3e3: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_f73614f348: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_3763fd75ee: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x130,
      clk => clk_1_sg_x130,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x130,
      clk => clk_1_sg_x130,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_4c0b07c2d5: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x130,
      clk => clk_1_sg_x130,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_e43eb2f177: entity work.twiddle_entity_e43eb2f177
    port map (
      ai => delay_q_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x130,
      clk_1 => clk_1_sg_x130,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/delay_b"

entity delay_b_entity_2f446d46db is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_2f446d46db;

architecture structural of delay_b_entity_2f446d46db is
  signal ce_1_sg_x131: std_logic;
  signal clk_1_sg_x131: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x131 <= ce_1;
  clk_1_sg_x131 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= delay_q_net_x3;

  delay: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x131,
      clk => clk_1_sg_x131,
      clr => '0',
      d => mux1_y_net_x0,
      q => delay_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11/sync_delay"

entity sync_delay_entity_1bb127f633 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_1bb127f633;

architecture structural of sync_delay_entity_1bb127f633 is
  signal ce_1_sg_x133: std_logic;
  signal clk_1_sg_x133: std_logic;
  signal constant1_op_net: std_logic_vector(2 downto 0);
  signal constant2_op_net: std_logic_vector(2 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(2 downto 0);
  signal counter_op_net: std_logic_vector(2 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x133 <= ce_1;
  clk_1_sg_x133 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a1c496ea88
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_3a3ea2f70b8548a5",
      op_arith => xlUnsigned,
      op_width => 3
    )
    port map (
      ce => ce_1_sg_x133,
      clk => clk_1_sg_x133,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_8fc7f5539b
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_47b317dab6
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_11"

entity fft_stage_11_entity_4f6b9006ee is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_11_entity_4f6b9006ee;

architecture structural of fft_stage_11_entity_4f6b9006ee is
  signal ce_1_sg_x134: std_logic;
  signal clk_1_sg_x134: std_logic;
  signal counter_op_net: std_logic_vector(2 downto 0);
  signal delay0_q_net_x3: std_logic;
  signal delay0_q_net_x4: std_logic;
  signal delay_q_net_x0: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal delay_q_net_x4: std_logic_vector(35 downto 0);
  signal fft_shift_net_x2: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x134 <= ce_1;
  clk_1_sg_x134 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x14 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x2 <= shift;
  delay0_q_net_x3 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x15;
  sync_out <= delay0_q_net_x4;

  butterfly_direct_6a735ce8e8: entity work.butterfly_direct_entity_6a735ce8e8
    port map (
      a => delay_q_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x134,
      clk_1 => clk_1_sg_x134,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x15,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x4
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_efa60dbe2ed9d35a",
      op_arith => xlUnsigned,
      op_width => 3
    )
    port map (
      ce => ce_1_sg_x134,
      clk => clk_1_sg_x134,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x3,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x134,
      clk => clk_1_sg_x134,
      clr => '0',
      d(0) => delay0_q_net_x3,
      q(0) => delay_q_net_x0
    );

  delay_b_2f446d46db: entity work.delay_b_entity_2f446d46db
    port map (
      ce_1 => ce_1_sg_x134,
      clk_1 => clk_1_sg_x134,
      din => mux1_y_net_x0,
      dout => delay_q_net_x3
    );

  delay_f_876cbfbaae: entity work.delay_b_entity_2f446d46db
    port map (
      ce_1 => ce_1_sg_x134,
      clk_1 => clk_1_sg_x134,
      din => reinterpret1_output_port_net_x14,
      dout => delay_q_net_x4
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x134,
      clk => clk_1_sg_x134,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x134,
      clk => clk_1_sg_x134,
      clr => '0',
      d0 => delay_q_net_x4,
      d1 => reinterpret2_output_port_net_x3,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x134,
      clk => clk_1_sg_x134,
      clr => '0',
      d0 => reinterpret2_output_port_net_x3,
      d1 => delay_q_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x2,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_1bb127f633: entity work.sync_delay_entity_1bb127f633
    port map (
      ce_1 => ce_1_sg_x134,
      clk_1 => clk_1_sg_x134,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_4ce9346ae0 is
  port (
    in_x0: in std_logic_vector(10 downto 0); 
    out_x0: out std_logic_vector(10 downto 0)
  );
end bit_reverse_entity_4ce9346ae0;

architecture structural of bit_reverse_entity_4ce9346ae0 is
  signal bit0_y_net: std_logic;
  signal bit10_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(10 downto 0);
  signal slice_y_net_x0: std_logic_vector(10 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit10: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit10_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_a0fa71d0d3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in10(0) => bit10_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_2f5130c631 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(10 downto 0); 
    add: out std_logic_vector(10 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_2f5130c631;

architecture structural of add_convert0_entity_2f5130c631 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(10 downto 0);
  signal ce_1_sg_x161: std_logic;
  signal clk_1_sg_x161: std_logic;
  signal concat_y_net: std_logic_vector(11 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal delay13_q_net: std_logic_vector(10 downto 0);
  signal delay14_q_net: std_logic_vector(10 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(11 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(9 downto 0);
  signal new_add_y_net: std_logic_vector(10 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x161 <= ce_1;
  clk_1_sg_x161 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_7ad1e33701
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 11,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 11,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9769d05421
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 12,
      y_width => 11
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_0d93032837 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(10 downto 0); 
    add: out std_logic_vector(10 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_0d93032837;

architecture structural of add_convert1_entity_0d93032837 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(10 downto 0);
  signal ce_1_sg_x162: std_logic;
  signal clk_1_sg_x162: std_logic;
  signal concat_y_net: std_logic_vector(11 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal delay13_q_net: std_logic_vector(10 downto 0);
  signal delay14_q_net: std_logic_vector(10 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(11 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(9 downto 0);
  signal new_add_y_net: std_logic_vector(10 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x162 <= ce_1;
  clk_1_sg_x162 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_7ad1e33701
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 11,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 11,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x162,
      clk => clk_1_sg_x162,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9769d05421
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 12,
      y_width => 11
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_6eb639ceaa is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(10 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_6eb639ceaa;

architecture structural of cosin_entity_6eb639ceaa is
  signal assert_dout_net_x1: std_logic_vector(10 downto 0);
  signal ce_1_sg_x165: std_logic;
  signal clk_1_sg_x165: std_logic;
  signal concat_y_net_x1: std_logic_vector(10 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(10 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x165 <= ce_1;
  clk_1_sg_x165 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_2f5130c631: entity work.add_convert0_entity_2f5130c631
    port map (
      ce_1 => ce_1_sg_x165,
      clk_1 => clk_1_sg_x165,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_0d93032837: entity work.add_convert1_entity_0d93032837
    port map (
      ce_1 => ce_1_sg_x165,
      clk_1 => clk_1_sg_x165,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 11,
      dout_width => 11
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x165,
      clk => clk_1_sg_x165,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x165,
      clk => clk_1_sg_x165,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x165,
      clk => clk_1_sg_x165,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_c4175667d0: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x165,
      clk_1 => clk_1_sg_x165,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_1956ff7d54: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x165,
      clk_1 => clk_1_sg_x165,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_core
    generic map (
      c_address_width_a => 11,
      c_address_width_b => 11,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_488bc588e4c66edf",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x165,
      a_clk => clk_1_sg_x165,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x165,
      b_clk => clk_1_sg_x165,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_5eba3a6b84 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_5eba3a6b84;

architecture structural of coeff_gen_entity_5eba3a6b84 is
  signal ce_1_sg_x166: std_logic;
  signal clk_1_sg_x166: std_logic;
  signal concat_y_net_x1: std_logic_vector(10 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(10 downto 0);

begin
  ce_1_sg_x166 <= ce_1;
  clk_1_sg_x166 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_4ce9346ae0: entity work.bit_reverse_entity_4ce9346ae0
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_6eb639ceaa: entity work.cosin_entity_6eb639ceaa
    port map (
      ce_1 => ce_1_sg_x166,
      clk_1 => clk_1_sg_x166,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x166,
      clk => clk_1_sg_x166,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_ac34020bca: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 11,
      x_width => 12,
      y_width => 11
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct/twiddle"

entity twiddle_entity_33ed0ffacc is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_33ed0ffacc;

architecture structural of twiddle_entity_33ed0ffacc is
  signal ce_1_sg_x167: std_logic;
  signal clk_1_sg_x167: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal delay_q_net_x1: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  delay_q_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x167 <= ce_1;
  clk_1_sg_x167 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_82e00ff98b: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x167,
      clk_1 => clk_1_sg_x167,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_ba93af5cc8: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => delay_q_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_99b4f46432: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_af3f352a8a: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_4bb10f5c74: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x167,
      clk_1 => clk_1_sg_x167,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_5eba3a6b84: entity work.coeff_gen_entity_5eba3a6b84
    port map (
      ce_1 => ce_1_sg_x167,
      clk_1 => clk_1_sg_x167,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/butterfly_direct"

entity butterfly_direct_entity_d133aef3f3 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_d133aef3f3;

architecture structural of butterfly_direct_entity_d133aef3f3 is
  signal ce_1_sg_x168: std_logic;
  signal clk_1_sg_x168: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal delay_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  delay_q_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x168 <= ce_1;
  clk_1_sg_x168 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_2a88d8383a: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      dout => concatenate_y_net_x3
    );

  bus_convert_c48bfbae81: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_4d2fe298c2: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_ce245c83ba: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_403e21fa27: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_12c24e83ce: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_fb8107f421: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_1361386295: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x168,
      clk => clk_1_sg_x168,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x168,
      clk => clk_1_sg_x168,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_f567a9b0ee: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x168,
      clk => clk_1_sg_x168,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_33ed0ffacc: entity work.twiddle_entity_33ed0ffacc
    port map (
      ai => delay_q_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x168,
      clk_1 => clk_1_sg_x168,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/delay_b"

entity delay_b_entity_2438f8654b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_2438f8654b;

architecture structural of delay_b_entity_2438f8654b is
  signal ce_1_sg_x169: std_logic;
  signal clk_1_sg_x169: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x169 <= ce_1;
  clk_1_sg_x169 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= delay_q_net_x3;

  delay: entity work.delay_38898c80c0
    port map (
      ce => ce_1_sg_x169,
      clk => clk_1_sg_x169,
      clr => '0',
      d => mux1_y_net_x0,
      q => delay_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12/sync_delay"

entity sync_delay_entity_ba1ce49596 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_ba1ce49596;

architecture structural of sync_delay_entity_ba1ce49596 is
  signal ce_1_sg_x171: std_logic;
  signal clk_1_sg_x171: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x171 <= ce_1;
  clk_1_sg_x171 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_99383d874600f8be",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x171,
      clk => clk_1_sg_x171,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f9928864ea
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_12"

entity fft_stage_12_entity_4d66daf6cf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_12_entity_4d66daf6cf;

architecture structural of fft_stage_12_entity_4d66daf6cf is
  signal ce_1_sg_x172: std_logic;
  signal clk_1_sg_x172: std_logic;
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay_q_net_x0: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal delay_q_net_x4: std_logic_vector(35 downto 0);
  signal fft_shift_net_x3: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x172 <= ce_1;
  clk_1_sg_x172 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x17 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x3 <= shift;
  delay0_q_net_x5 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x12;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_d133aef3f3: entity work.butterfly_direct_entity_d133aef3f3
    port map (
      a => delay_q_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x172,
      clk_1 => clk_1_sg_x172,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x12,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_533dcbdd307dbf50",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x172,
      clk => clk_1_sg_x172,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x5,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x172,
      clk => clk_1_sg_x172,
      clr => '0',
      d(0) => delay0_q_net_x5,
      q(0) => delay_q_net_x0
    );

  delay_b_2438f8654b: entity work.delay_b_entity_2438f8654b
    port map (
      ce_1 => ce_1_sg_x172,
      clk_1 => clk_1_sg_x172,
      din => mux1_y_net_x0,
      dout => delay_q_net_x3
    );

  delay_f_33d5a77eca: entity work.delay_b_entity_2438f8654b
    port map (
      ce_1 => ce_1_sg_x172,
      clk_1 => clk_1_sg_x172,
      din => reinterpret1_output_port_net_x17,
      dout => delay_q_net_x4
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x172,
      clk => clk_1_sg_x172,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x172,
      clk => clk_1_sg_x172,
      clr => '0',
      d0 => delay_q_net_x4,
      d1 => reinterpret2_output_port_net_x5,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x172,
      clk => clk_1_sg_x172,
      clr => '0',
      d0 => reinterpret2_output_port_net_x5,
      d1 => delay_q_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x3,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_ba1ce49596: entity work.sync_delay_entity_ba1ce49596
    port map (
      ce_1 => ce_1_sg_x172,
      clk_1 => clk_1_sg_x172,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_a889b2a85c is
  port (
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(11 downto 0)
  );
end bit_reverse_entity_a889b2a85c;

architecture structural of bit_reverse_entity_a889b2a85c is
  signal bit0_y_net: std_logic;
  signal bit10_y_net: std_logic;
  signal bit11_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(11 downto 0);
  signal slice_y_net_x0: std_logic_vector(11 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit10: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit10_y_net
    );

  bit11: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit11_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_ef66525e56
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in10(0) => bit10_y_net,
      in11(0) => bit11_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_6e803c8dba is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(11 downto 0); 
    add: out std_logic_vector(11 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_6e803c8dba;

architecture structural of add_convert0_entity_6e803c8dba is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(11 downto 0);
  signal ce_1_sg_x199: std_logic;
  signal clk_1_sg_x199: std_logic;
  signal concat_y_net: std_logic_vector(12 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(11 downto 0);
  signal delay13_q_net: std_logic_vector(11 downto 0);
  signal delay14_q_net: std_logic_vector(11 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(12 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(10 downto 0);
  signal new_add_y_net: std_logic_vector(11 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x199 <= ce_1;
  clk_1_sg_x199 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_8503582fb5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 12,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 12,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_118109a960
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 12,
      x_width => 13,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_22344e2a75 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(11 downto 0); 
    add: out std_logic_vector(11 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_22344e2a75;

architecture structural of add_convert1_entity_22344e2a75 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(11 downto 0);
  signal ce_1_sg_x200: std_logic;
  signal clk_1_sg_x200: std_logic;
  signal concat_y_net: std_logic_vector(12 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(11 downto 0);
  signal delay13_q_net: std_logic_vector(11 downto 0);
  signal delay14_q_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(12 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(10 downto 0);
  signal new_add_y_net: std_logic_vector(11 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x200 <= ce_1;
  clk_1_sg_x200 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_8503582fb5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 12,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 12,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x200,
      clk => clk_1_sg_x200,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_118109a960
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 12,
      x_width => 13,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_4f13fc5a71 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(11 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_4f13fc5a71;

architecture structural of cosin_entity_4f13fc5a71 is
  signal assert_dout_net_x1: std_logic_vector(11 downto 0);
  signal ce_1_sg_x203: std_logic;
  signal clk_1_sg_x203: std_logic;
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(11 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(11 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x203 <= ce_1;
  clk_1_sg_x203 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_6e803c8dba: entity work.add_convert0_entity_6e803c8dba
    port map (
      ce_1 => ce_1_sg_x203,
      clk_1 => clk_1_sg_x203,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_22344e2a75: entity work.add_convert1_entity_22344e2a75
    port map (
      ce_1 => ce_1_sg_x203,
      clk_1 => clk_1_sg_x203,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 12,
      dout_width => 12
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x203,
      clk => clk_1_sg_x203,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x203,
      clk => clk_1_sg_x203,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x203,
      clk => clk_1_sg_x203,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_6c850d0e45: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x203,
      clk_1 => clk_1_sg_x203,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_e468a3ac30: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x203,
      clk_1 => clk_1_sg_x203,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_core
    generic map (
      c_address_width_a => 12,
      c_address_width_b => 12,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_53d3a85261e207bb",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x203,
      a_clk => clk_1_sg_x203,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x203,
      b_clk => clk_1_sg_x203,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_552fac7a8c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_552fac7a8c;

architecture structural of coeff_gen_entity_552fac7a8c is
  signal ce_1_sg_x204: std_logic;
  signal clk_1_sg_x204: std_logic;
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x204 <= ce_1;
  clk_1_sg_x204 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_a889b2a85c: entity work.bit_reverse_entity_a889b2a85c
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_4f13fc5a71: entity work.cosin_entity_4f13fc5a71
    port map (
      ce_1 => ce_1_sg_x204,
      clk_1 => clk_1_sg_x204,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x204,
      clk => clk_1_sg_x204,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_23e8c8bac6: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 12,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct/twiddle"

entity twiddle_entity_75a6f99351 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_75a6f99351;

architecture structural of twiddle_entity_75a6f99351 is
  signal ce_1_sg_x205: std_logic;
  signal clk_1_sg_x205: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal delay_q_net_x1: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  delay_q_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x205 <= ce_1;
  clk_1_sg_x205 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_dc956d4b82: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x205,
      clk_1 => clk_1_sg_x205,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_900907d88b: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => delay_q_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_e0344067c0: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_7b8f10b1c0: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_8ef43c2602: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x205,
      clk_1 => clk_1_sg_x205,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_552fac7a8c: entity work.coeff_gen_entity_552fac7a8c
    port map (
      ce_1 => ce_1_sg_x205,
      clk_1 => clk_1_sg_x205,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/butterfly_direct"

entity butterfly_direct_entity_f7d3b38784 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_f7d3b38784;

architecture structural of butterfly_direct_entity_f7d3b38784 is
  signal ce_1_sg_x206: std_logic;
  signal clk_1_sg_x206: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x3: std_logic;
  signal delay2_q_net: std_logic;
  signal delay_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  delay_q_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x206 <= ce_1;
  clk_1_sg_x206 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x3;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x3;

  bus_add_3ac32c4378: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      dout => concatenate_y_net_x3
    );

  bus_convert_e0cb53f184: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_e89cea9f62: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_norm0_be5f445594: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_b018d4e3d1: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_75685eb826: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_7ab0f1679b: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_75d205b5b9: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x206,
      clk => clk_1_sg_x206,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x3
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x206,
      clk => clk_1_sg_x206,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_ad161f32ec: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x206,
      clk => clk_1_sg_x206,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_75a6f99351: entity work.twiddle_entity_75a6f99351
    port map (
      ai => delay_q_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x206,
      clk_1 => clk_1_sg_x206,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/delay_b"

entity delay_b_entity_198843ae55 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_198843ae55;

architecture structural of delay_b_entity_198843ae55 is
  signal ce_1_sg_x207: std_logic;
  signal clk_1_sg_x207: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x207 <= ce_1;
  clk_1_sg_x207 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= delay_q_net_x3;

  delay: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x207,
      clk => clk_1_sg_x207,
      clr => '0',
      d => mux1_y_net_x0,
      q => delay_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13/sync_delay"

entity sync_delay_entity_a89ef53aef is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_a89ef53aef;

architecture structural of sync_delay_entity_a89ef53aef is
  signal ce_1_sg_x209: std_logic;
  signal clk_1_sg_x209: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x209 <= ce_1;
  clk_1_sg_x209 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_99383d874600f8be",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x209,
      clk => clk_1_sg_x209,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f9928864ea
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_13"

entity fft_stage_13_entity_02afd91842 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_13_entity_02afd91842;

architecture structural of fft_stage_13_entity_02afd91842 is
  signal ce_1_sg_x210: std_logic;
  signal clk_1_sg_x210: std_logic;
  signal counter_op_net: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x4: std_logic;
  signal delay_q_net_x0: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal delay_q_net_x4: std_logic_vector(35 downto 0);
  signal fft_shift_net_x4: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x8: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x210 <= ce_1;
  clk_1_sg_x210 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x14 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x4 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x8;
  out2 <= reinterpret1_output_port_net_x15;
  sync_out <= delay0_q_net_x4;

  butterfly_direct_f7d3b38784: entity work.butterfly_direct_entity_f7d3b38784
    port map (
      a => delay_q_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x210,
      clk_1 => clk_1_sg_x210,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x15,
      a_bw_x0 => reinterpret2_output_port_net_x8,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x4
    );

  counter: entity work.counter_9b03e3d644
    port map (
      ce => ce_1_sg_x210,
      clk => clk_1_sg_x210,
      clr => '0',
      rst(0) => delay0_q_net_x2,
      op(0) => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x210,
      clk => clk_1_sg_x210,
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => delay_q_net_x0
    );

  delay_b_198843ae55: entity work.delay_b_entity_198843ae55
    port map (
      ce_1 => ce_1_sg_x210,
      clk_1 => clk_1_sg_x210,
      din => mux1_y_net_x0,
      dout => delay_q_net_x3
    );

  delay_f_a103f8b8fe: entity work.delay_b_entity_198843ae55
    port map (
      ce_1 => ce_1_sg_x210,
      clk_1 => clk_1_sg_x210,
      din => reinterpret1_output_port_net_x14,
      dout => delay_q_net_x4
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x210,
      clk => clk_1_sg_x210,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x210,
      clk => clk_1_sg_x210,
      clr => '0',
      d0 => delay_q_net_x4,
      d1 => reinterpret2_output_port_net_x7,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x210,
      clk => clk_1_sg_x210,
      clr => '0',
      d0 => reinterpret2_output_port_net_x7,
      d1 => delay_q_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x4,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 1,
      y_width => 1
    )
    port map (
      x(0) => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_a89ef53aef: entity work.sync_delay_entity_a89ef53aef
    port map (
      ce_1 => ce_1_sg_x210,
      clk_1 => clk_1_sg_x210,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2/butterfly_direct/twiddle/negate"

entity negate_entity_90afb2f493 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(17 downto 0); 
    dout: out std_logic_vector(17 downto 0)
  );
end negate_entity_90afb2f493;

architecture structural of negate_entity_90afb2f493 is
  signal ce_1_sg_x228: std_logic;
  signal clk_1_sg_x228: std_logic;
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x228 <= ce_1;
  clk_1_sg_x228 <= clk_1;
  reinterpret2_output_port_net_x2 <= din;
  dout <= reinterpret1_output_port_net_x2;

  bussify_4c1a10b553: entity work.bussify_entity_427b04c969
    port map (
      in1 => neg1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

  debus_3c23ef0562: entity work.a_debus_entity_459b56afaf
    port map (
      bus_in => reinterpret2_output_port_net_x2,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  neg1: entity work.negate_894f23b88c
    port map (
      ce => ce_1_sg_x228,
      clk => clk_1_sg_x228,
      clr => '0',
      ip => reinterpret1_output_port_net_x1,
      op => neg1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2/butterfly_direct/twiddle"

entity twiddle_entity_379d88ebbf is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_379d88ebbf;

architecture structural of twiddle_entity_379d88ebbf is
  signal ce_1_sg_x229: std_logic;
  signal clk_1_sg_x229: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay0_q_net_x4: std_logic_vector(35 downto 0);
  signal delay2_q_net: std_logic;
  signal delay3_q_net: std_logic_vector(17 downto 0);
  signal delay4_q_net: std_logic_vector(17 downto 0);
  signal delay5_q_net: std_logic_vector(17 downto 0);
  signal delay6_q_net: std_logic_vector(17 downto 0);
  signal delay7_q_net: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal mux0_y_net_x0: std_logic_vector(17 downto 0);
  signal mux1_y_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal slice_y_net: std_logic;

begin
  ram_data_out_net_x0 <= ai;
  mux_y_net_x1 <= bi;
  ce_1_sg_x229 <= ce_1;
  clk_1_sg_x229 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= delay0_q_net_x4;
  bwo <= reinterpret_out_output_port_net_x5;
  sync_out <= delay8_q_net_x0;

  bus_create_5286d58582: entity work.join_entity_dce4ac7e98
    port map (
      in1 => mux0_y_net_x0,
      in2 => mux1_y_net_x0,
      bus_out => concatenate_y_net_x2
    );

  bus_expand_5fb439edb0: entity work.bus_expand_a_entity_e0cf78c6cc
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x2
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      rst(0) => delay7_q_net,
      op => counter_op_net
    );

  delay0: entity work.delay_4c85700954
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => ram_data_out_net_x0,
      q => delay0_q_net_x4
    );

  delay2: entity work.delay_5b3ce5f2ae
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d(0) => slice_y_net,
      q(0) => delay2_q_net
    );

  delay3: entity work.delay_4217913c13
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => delay6_q_net,
      q => delay3_q_net
    );

  delay4: entity work.delay_c462a80bee
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => reinterpret1_output_port_net_x2,
      q => delay4_q_net
    );

  delay5: entity work.delay_328e8ebbb5
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => reinterpret2_output_port_net_x2,
      q => delay5_q_net
    );

  delay6: entity work.delay_328e8ebbb5
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => delay6_q_net
    );

  delay7: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d(0) => mux_y_net_x2,
      q(0) => delay7_q_net
    );

  delay8: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d(0) => delay7_q_net,
      q(0) => delay8_q_net_x0
    );

  munge_in_6211aa3173: entity work.munge_a_entity_40c03aaddb
    port map (
      din => mux_y_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_out_5e592e090a: entity work.munge_a_entity_40c03aaddb
    port map (
      din => concatenate_y_net_x2,
      dout => reinterpret_out_output_port_net_x5
    );

  mux0: entity work.mux_30e9ca90db
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d0 => delay5_q_net,
      d1 => delay6_q_net,
      sel(0) => slice_y_net,
      y => mux0_y_net_x0
    );

  mux1: entity work.mux_181e58d842
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d0 => delay3_q_net,
      d1 => delay4_q_net,
      sel(0) => delay2_q_net,
      y => mux1_y_net_x0
    );

  negate_90afb2f493: entity work.negate_entity_90afb2f493
    port map (
      ce_1 => ce_1_sg_x229,
      clk_1 => clk_1_sg_x229,
      din => reinterpret2_output_port_net_x2,
      dout => reinterpret1_output_port_net_x2
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2/butterfly_direct"

entity butterfly_direct_entity_e7cfb99339 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_e7cfb99339;

architecture structural of butterfly_direct_entity_e7cfb99339 is
  signal ce_1_sg_x230: std_logic;
  signal clk_1_sg_x230: std_logic;
  signal concat_y_net_x3: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay0_q_net_x4: std_logic_vector(35 downto 0);
  signal delay2_q_net: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal mux_y_net_x2: std_logic_vector(79 downto 0);
  signal mux_y_net_x4: std_logic_vector(35 downto 0);
  signal mux_y_net_x5: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x1 <= a;
  mux_y_net_x4 <= b;
  ce_1_sg_x230 <= ce_1;
  clk_1_sg_x230 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x5 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x5;
  sync_out <= delay0_q_net_x0;

  bus_add_3d0e740a18: entity work.bus_add_entity_695cb26b69
    port map (
      a => delay0_q_net_x4,
      b => reinterpret_out_output_port_net_x5,
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      dout => concatenate_y_net_x1
    );

  bus_convert_9164ba6aff: entity work.bus_convert_entity_82369b5cdf
    port map (
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      din => mux_y_net_x2,
      dout => concatenate_y_net_x3,
      overflow => concatenate_y_net_x4
    );

  bus_expand_4778bf4ba8: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_1adca9e1e9: entity work.bus_norm0_entity_f70daa5f43
    port map (
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x5
    );

  bus_norm1_56535b5a2c: entity work.bus_norm1_entity_1de1ca87af
    port map (
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_eb1b3be6fb: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x5
    );

  bus_scale_b4b6296b21: entity work.bus_scale_entity_472dd14792
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_109da66520: entity work.bus_sub_entity_2925aed405
    port map (
      a => delay0_q_net_x4,
      b => reinterpret_out_output_port_net_x5,
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_4822199898
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x1,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d(0) => delay8_q_net_x0,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_aafba4c121: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x4,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_9ff8aec2dc
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d0 => concatenate_y_net_x5,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x2
    );

  twiddle_379d88ebbf: entity work.twiddle_entity_379d88ebbf
    port map (
      ai => ram_data_out_net_x1,
      bi => mux_y_net_x4,
      ce_1 => ce_1_sg_x230,
      clk_1 => clk_1_sg_x230,
      sync_in => mux_y_net_x5,
      ao => delay0_q_net_x4,
      bwo => reinterpret_out_output_port_net_x5,
      sync_out => delay8_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2/delay_b"

entity delay_b_entity_a5401bb008 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_a5401bb008;

architecture structural of delay_b_entity_a5401bb008 is
  signal ce_1_sg_x231: std_logic;
  signal clk_1_sg_x231: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(10 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x231 <= ce_1;
  clk_1_sg_x231 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x2;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 2044,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_60602034a1d84a16",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 11
    )
    port map (
      ce => ce_1_sg_x231,
      clk => clk_1_sg_x231,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 11,
      c_width => 36,
      core_name0 => "bmg_72_7e8fa68244af6cff",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x231,
      clk => clk_1_sg_x231,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2/sync_delay"

entity sync_delay_entity_9ee9307058 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_9ee9307058;

architecture structural of sync_delay_entity_9ee9307058 is
  signal ce_1_sg_x233: std_logic;
  signal clk_1_sg_x233: std_logic;
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(11 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x6: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x233 <= ce_1;
  clk_1_sg_x233 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x6;

  constant1: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_7c91b1b314
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_a2916e7e77833dd6",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x233,
      clk => clk_1_sg_x233,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x6
    );

  relational: entity work.relational_d36fe12c1c
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_acb3c05dd0
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_2"

entity fft_stage_2_entity_012e00c14b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_2_entity_012e00c14b;

architecture structural of fft_stage_2_entity_012e00c14b is
  signal ce_1_sg_x234: std_logic;
  signal clk_1_sg_x234: std_logic;
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x5: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic_vector(35 downto 0);
  signal mux_y_net_x6: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x234 <= ce_1;
  clk_1_sg_x234 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x8 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x5 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x9;
  sync_out <= delay0_q_net_x3;

  butterfly_direct_e7cfb99339: entity work.butterfly_direct_entity_e7cfb99339
    port map (
      a => ram_data_out_net_x2,
      b => mux_y_net_x4,
      ce_1 => ce_1_sg_x234,
      clk_1 => clk_1_sg_x234,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x6,
      a_bw => reinterpret1_output_port_net_x9,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x5,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x2,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => delay_q_net_x0
    );

  delay_b_a5401bb008: entity work.delay_b_entity_a5401bb008
    port map (
      ce_1 => ce_1_sg_x234,
      clk_1 => clk_1_sg_x234,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x2
    );

  delay_f_5a950dbeff: entity work.delay_b_entity_a5401bb008
    port map (
      ce_1 => ce_1_sg_x234,
      clk_1 => clk_1_sg_x234,
      din => reinterpret1_output_port_net_x8,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x5,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x3,
      sel(0) => slice1_y_net,
      y => mux_y_net_x4
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      d0 => reinterpret2_output_port_net_x3,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x5,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_9ee9307058: entity work.sync_delay_entity_9ee9307058
    port map (
      ce_1 => ce_1_sg_x234,
      clk_1 => clk_1_sg_x234,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x6
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_b4fce180d8 is
  port (
    in_x0: in std_logic_vector(1 downto 0); 
    out_x0: out std_logic_vector(1 downto 0)
  );
end bit_reverse_entity_b4fce180d8;

architecture structural of bit_reverse_entity_b4fce180d8 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(1 downto 0);
  signal slice_y_net_x0: std_logic_vector(1 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  concat: entity work.concat_e6f5ee726b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_dc18c9584e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(1 downto 0); 
    add: out std_logic_vector(1 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_dc18c9584e;

architecture structural of add_convert0_entity_dc18c9584e is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(1 downto 0);
  signal ce_1_sg_x261: std_logic;
  signal clk_1_sg_x261: std_logic;
  signal concat_y_net: std_logic_vector(2 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal delay13_q_net: std_logic_vector(1 downto 0);
  signal delay14_q_net: std_logic_vector(1 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(2 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic;
  signal new_add_y_net: std_logic_vector(1 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x261 <= ce_1;
  clk_1_sg_x261 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_6160d7387c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1(0) => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 2,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 2,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_4a9a9a25a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => fluff_y_net,
      y(0) => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 2,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_d76a56f639 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(1 downto 0); 
    add: out std_logic_vector(1 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_d76a56f639;

architecture structural of add_convert1_entity_d76a56f639 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(1 downto 0);
  signal ce_1_sg_x262: std_logic;
  signal clk_1_sg_x262: std_logic;
  signal concat_y_net: std_logic_vector(2 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal delay13_q_net: std_logic_vector(1 downto 0);
  signal delay14_q_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(2 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic;
  signal new_add_y_net: std_logic_vector(1 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x262 <= ce_1;
  clk_1_sg_x262 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_6160d7387c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1(0) => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 2,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 2,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_4a9a9a25a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => fluff_y_net,
      y(0) => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 2,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_68c0ea6425 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(1 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_68c0ea6425;

architecture structural of cosin_entity_68c0ea6425 is
  signal assert_dout_net_x1: std_logic_vector(1 downto 0);
  signal ce_1_sg_x265: std_logic;
  signal clk_1_sg_x265: std_logic;
  signal concat_y_net_x1: std_logic_vector(1 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(1 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x265 <= ce_1;
  clk_1_sg_x265 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_dc18c9584e: entity work.add_convert0_entity_dc18c9584e
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_d76a56f639: entity work.add_convert1_entity_d76a56f639
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 2,
      dout_width => 2
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_3d81cbdfe4: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_16d2db8745: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_core
    generic map (
      addr_width => 2,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_505931c5b3ea228e",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x265,
      a_clk => clk_1_sg_x265,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x265,
      b_clk => clk_1_sg_x265,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_ad3a81b5c0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_ad3a81b5c0;

architecture structural of coeff_gen_entity_ad3a81b5c0 is
  signal ce_1_sg_x266: std_logic;
  signal clk_1_sg_x266: std_logic;
  signal concat_y_net_x1: std_logic_vector(1 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x266 <= ce_1;
  clk_1_sg_x266 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_b4fce180d8: entity work.bit_reverse_entity_b4fce180d8
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_68c0ea6425: entity work.cosin_entity_68c0ea6425
    port map (
      ce_1 => ce_1_sg_x266,
      clk_1 => clk_1_sg_x266,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x266,
      clk => clk_1_sg_x266,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_495ae8a001: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct/twiddle"

entity twiddle_entity_b90d438adc is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_b90d438adc;

architecture structural of twiddle_entity_b90d438adc is
  signal ce_1_sg_x267: std_logic;
  signal clk_1_sg_x267: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x267 <= ce_1;
  clk_1_sg_x267 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_33f279bae1: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x267,
      clk_1 => clk_1_sg_x267,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_64225822e4: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_2c42e8fd1e: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_7e4d9192ed: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_4bbd37883a: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x267,
      clk_1 => clk_1_sg_x267,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_ad3a81b5c0: entity work.coeff_gen_entity_ad3a81b5c0
    port map (
      ce_1 => ce_1_sg_x267,
      clk_1 => clk_1_sg_x267,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/butterfly_direct"

entity butterfly_direct_entity_e0e9981582 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_e0e9981582;

architecture structural of butterfly_direct_entity_e0e9981582 is
  signal ce_1_sg_x268: std_logic;
  signal clk_1_sg_x268: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x268 <= ce_1;
  clk_1_sg_x268 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_341faea5ce: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      dout => concatenate_y_net_x3
    );

  bus_convert_eea6f1b583: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_ae88b2b997: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_b6cfbb11fb: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_6da21410a4: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_96bb02e1e5: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_c83199e3d7: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_f1636466ab: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x268,
      clk => clk_1_sg_x268,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x268,
      clk => clk_1_sg_x268,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_9c76c4f36b: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x268,
      clk => clk_1_sg_x268,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_b90d438adc: entity work.twiddle_entity_b90d438adc
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x268,
      clk_1 => clk_1_sg_x268,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/delay_b"

entity delay_b_entity_a58de5738f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_a58de5738f;

architecture structural of delay_b_entity_a58de5738f is
  signal ce_1_sg_x269: std_logic;
  signal clk_1_sg_x269: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x269 <= ce_1;
  clk_1_sg_x269 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 1020,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_89850cbcf0fde6e9",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x269,
      clk => clk_1_sg_x269,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 10,
      c_width => 36,
      core_name0 => "bmg_72_756e5f183b33a31a",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x269,
      clk => clk_1_sg_x269,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3/sync_delay"

entity sync_delay_entity_3dadc1273e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_3dadc1273e;

architecture structural of sync_delay_entity_3dadc1273e is
  signal ce_1_sg_x271: std_logic;
  signal clk_1_sg_x271: std_logic;
  signal constant1_op_net: std_logic_vector(10 downto 0);
  signal constant2_op_net: std_logic_vector(10 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(10 downto 0);
  signal counter_op_net: std_logic_vector(10 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x271 <= ce_1;
  clk_1_sg_x271 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_a3923dd146
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_0604807f72
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_118598964d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_2f7113c203379501",
      op_arith => xlUnsigned,
      op_width => 11
    )
    port map (
      ce => ce_1_sg_x271,
      clk => clk_1_sg_x271,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_2147430058
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_b4b277ae0f
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_3"

entity fft_stage_3_entity_33ea5e4989 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_3_entity_33ea5e4989;

architecture structural of fft_stage_3_entity_33ea5e4989 is
  signal ce_1_sg_x272: std_logic;
  signal clk_1_sg_x272: std_logic;
  signal counter_op_net: std_logic_vector(10 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x6: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x272 <= ce_1;
  clk_1_sg_x272 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x12 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x6 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x13;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_e0e9981582: entity work.butterfly_direct_entity_e0e9981582
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x272,
      clk_1 => clk_1_sg_x272,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x13,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_60602034a1d84a16",
      op_arith => xlUnsigned,
      op_width => 11
    )
    port map (
      ce => ce_1_sg_x272,
      clk => clk_1_sg_x272,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x4,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x272,
      clk => clk_1_sg_x272,
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => delay_q_net_x0
    );

  delay_b_a58de5738f: entity work.delay_b_entity_a58de5738f
    port map (
      ce_1 => ce_1_sg_x272,
      clk_1 => clk_1_sg_x272,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_3d8cf3a7fb: entity work.delay_b_entity_a58de5738f
    port map (
      ce_1 => ce_1_sg_x272,
      clk_1 => clk_1_sg_x272,
      din => reinterpret1_output_port_net_x12,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x272,
      clk => clk_1_sg_x272,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x272,
      clk => clk_1_sg_x272,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x5,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x272,
      clk => clk_1_sg_x272,
      clr => '0',
      d0 => reinterpret2_output_port_net_x5,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x6,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_3dadc1273e: entity work.sync_delay_entity_3dadc1273e
    port map (
      ce_1 => ce_1_sg_x272,
      clk_1 => clk_1_sg_x272,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_e679e17e2b is
  port (
    in_x0: in std_logic_vector(2 downto 0); 
    out_x0: out std_logic_vector(2 downto 0)
  );
end bit_reverse_entity_e679e17e2b;

architecture structural of bit_reverse_entity_e679e17e2b is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(2 downto 0);
  signal slice_y_net_x0: std_logic_vector(2 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  concat: entity work.concat_452c4d3410
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_6a0feb5dcc is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(2 downto 0); 
    add: out std_logic_vector(2 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_6a0feb5dcc;

architecture structural of add_convert0_entity_6a0feb5dcc is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(2 downto 0);
  signal ce_1_sg_x299: std_logic;
  signal clk_1_sg_x299: std_logic;
  signal concat_y_net: std_logic_vector(3 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal delay13_q_net: std_logic_vector(2 downto 0);
  signal delay14_q_net: std_logic_vector(2 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(3 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(1 downto 0);
  signal new_add_y_net: std_logic_vector(2 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x299 <= ce_1;
  clk_1_sg_x299 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x299,
      clk => clk_1_sg_x299,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 3,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 3,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x299,
      clk => clk_1_sg_x299,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x299,
      clk => clk_1_sg_x299,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x299,
      clk => clk_1_sg_x299,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x299,
      clk => clk_1_sg_x299,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_949f038a6d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 4,
      y_width => 3
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_94be4a15f7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(2 downto 0); 
    add: out std_logic_vector(2 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_94be4a15f7;

architecture structural of add_convert1_entity_94be4a15f7 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(2 downto 0);
  signal ce_1_sg_x300: std_logic;
  signal clk_1_sg_x300: std_logic;
  signal concat_y_net: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal delay13_q_net: std_logic_vector(2 downto 0);
  signal delay14_q_net: std_logic_vector(2 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(3 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(1 downto 0);
  signal new_add_y_net: std_logic_vector(2 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x300 <= ce_1;
  clk_1_sg_x300 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 3,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 3,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x300,
      clk => clk_1_sg_x300,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_949f038a6d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 4,
      y_width => 3
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_bc43e3a4c5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(2 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_bc43e3a4c5;

architecture structural of cosin_entity_bc43e3a4c5 is
  signal assert_dout_net_x1: std_logic_vector(2 downto 0);
  signal ce_1_sg_x303: std_logic;
  signal clk_1_sg_x303: std_logic;
  signal concat_y_net_x1: std_logic_vector(2 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(2 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x303 <= ce_1;
  clk_1_sg_x303 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_6a0feb5dcc: entity work.add_convert0_entity_6a0feb5dcc
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_94be4a15f7: entity work.add_convert1_entity_94be4a15f7
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 3,
      dout_width => 3
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x303,
      clk => clk_1_sg_x303,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x303,
      clk => clk_1_sg_x303,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x303,
      clk => clk_1_sg_x303,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_e1fee0fd0d: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_7bcae090eb: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_core
    generic map (
      addr_width => 3,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_d20b02a9f8239c7a",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x303,
      a_clk => clk_1_sg_x303,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x303,
      b_clk => clk_1_sg_x303,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_d0f746b8cb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_d0f746b8cb;

architecture structural of coeff_gen_entity_d0f746b8cb is
  signal ce_1_sg_x304: std_logic;
  signal clk_1_sg_x304: std_logic;
  signal concat_y_net_x1: std_logic_vector(2 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(2 downto 0);

begin
  ce_1_sg_x304 <= ce_1;
  clk_1_sg_x304 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_e679e17e2b: entity work.bit_reverse_entity_e679e17e2b
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_bc43e3a4c5: entity work.cosin_entity_bc43e3a4c5
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x304,
      clk => clk_1_sg_x304,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_63189c15ea: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 11,
      x_width => 12,
      y_width => 3
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct/twiddle"

entity twiddle_entity_c5ce36f36f is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_c5ce36f36f;

architecture structural of twiddle_entity_c5ce36f36f is
  signal ce_1_sg_x305: std_logic;
  signal clk_1_sg_x305: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x305 <= ce_1;
  clk_1_sg_x305 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_a8597be60e: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x305,
      clk_1 => clk_1_sg_x305,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_32a9dee733: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_fe4e25d139: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_cd8554d55c: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_ddee2b7de1: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x305,
      clk_1 => clk_1_sg_x305,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_d0f746b8cb: entity work.coeff_gen_entity_d0f746b8cb
    port map (
      ce_1 => ce_1_sg_x305,
      clk_1 => clk_1_sg_x305,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/butterfly_direct"

entity butterfly_direct_entity_6ae06ea03e is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_6ae06ea03e;

architecture structural of butterfly_direct_entity_6ae06ea03e is
  signal ce_1_sg_x306: std_logic;
  signal clk_1_sg_x306: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x306 <= ce_1;
  clk_1_sg_x306 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_de8a533838: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      dout => concatenate_y_net_x3
    );

  bus_convert_c099a1336e: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_08b7316806: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_5b70207350: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_0c684f4a74: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_e8fe2e7a4e: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_0b58f086e3: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_2ea74fc977: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x306,
      clk => clk_1_sg_x306,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x306,
      clk => clk_1_sg_x306,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_de1e86bbf8: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x306,
      clk => clk_1_sg_x306,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_c5ce36f36f: entity work.twiddle_entity_c5ce36f36f
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x306,
      clk_1 => clk_1_sg_x306,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/delay_b"

entity delay_b_entity_e389d19113 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_e389d19113;

architecture structural of delay_b_entity_e389d19113 is
  signal ce_1_sg_x307: std_logic;
  signal clk_1_sg_x307: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x307 <= ce_1;
  clk_1_sg_x307 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 508,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_12b8e0a4a9ef4845",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x307,
      clk => clk_1_sg_x307,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 9,
      c_width => 36,
      core_name0 => "bmg_72_9fff5a02c6b3c277",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x307,
      clk => clk_1_sg_x307,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4/sync_delay"

entity sync_delay_entity_7ed60ac727 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_7ed60ac727;

architecture structural of sync_delay_entity_7ed60ac727 is
  signal ce_1_sg_x309: std_logic;
  signal clk_1_sg_x309: std_logic;
  signal constant1_op_net: std_logic_vector(9 downto 0);
  signal constant2_op_net: std_logic_vector(9 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(9 downto 0);
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x309 <= ce_1;
  clk_1_sg_x309 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_498bc68c14
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_fbc2f0cce1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_f1ac4bddff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_4adf855dd0e5af2a",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x309,
      clk => clk_1_sg_x309,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_0ffd72e037
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f6702ea2f7
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_4"

entity fft_stage_4_entity_a779b0edc3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_4_entity_a779b0edc3;

architecture structural of fft_stage_4_entity_a779b0edc3 is
  signal ce_1_sg_x310: std_logic;
  signal clk_1_sg_x310: std_logic;
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x7: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x310 <= ce_1;
  clk_1_sg_x310 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x15 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x7 <= shift;
  delay0_q_net_x6 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x16;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_6ae06ea03e: entity work.butterfly_direct_entity_6ae06ea03e
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x310,
      clk_1 => clk_1_sg_x310,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x16,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_89850cbcf0fde6e9",
      op_arith => xlUnsigned,
      op_width => 10
    )
    port map (
      ce => ce_1_sg_x310,
      clk => clk_1_sg_x310,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x6,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x310,
      clk => clk_1_sg_x310,
      clr => '0',
      d(0) => delay0_q_net_x6,
      q(0) => delay_q_net_x0
    );

  delay_b_e389d19113: entity work.delay_b_entity_e389d19113
    port map (
      ce_1 => ce_1_sg_x310,
      clk_1 => clk_1_sg_x310,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_400e03c913: entity work.delay_b_entity_e389d19113
    port map (
      ce_1 => ce_1_sg_x310,
      clk_1 => clk_1_sg_x310,
      din => reinterpret1_output_port_net_x15,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x310,
      clk => clk_1_sg_x310,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x310,
      clk => clk_1_sg_x310,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x7,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x310,
      clk => clk_1_sg_x310,
      clr => '0',
      d0 => reinterpret2_output_port_net_x7,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x7,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_7ed60ac727: entity work.sync_delay_entity_7ed60ac727
    port map (
      ce_1 => ce_1_sg_x310,
      clk_1 => clk_1_sg_x310,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_21d5d92029 is
  port (
    in_x0: in std_logic_vector(3 downto 0); 
    out_x0: out std_logic_vector(3 downto 0)
  );
end bit_reverse_entity_21d5d92029;

architecture structural of bit_reverse_entity_21d5d92029 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(3 downto 0);
  signal slice_y_net_x0: std_logic_vector(3 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  concat: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_a9a42ddd37 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(3 downto 0); 
    add: out std_logic_vector(3 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_a9a42ddd37;

architecture structural of add_convert0_entity_a9a42ddd37 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x337: std_logic;
  signal clk_1_sg_x337: std_logic;
  signal concat_y_net: std_logic_vector(4 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal delay13_q_net: std_logic_vector(3 downto 0);
  signal delay14_q_net: std_logic_vector(3 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(4 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(2 downto 0);
  signal new_add_y_net: std_logic_vector(3 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x337 <= ce_1;
  clk_1_sg_x337 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x337,
      clk => clk_1_sg_x337,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_8f12c32de0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 4,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 4,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x337,
      clk => clk_1_sg_x337,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x337,
      clk => clk_1_sg_x337,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x337,
      clk => clk_1_sg_x337,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x337,
      clk => clk_1_sg_x337,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_cf540617d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 5,
      y_width => 3
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 5,
      y_width => 4
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 5,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_50e644ef30 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(3 downto 0); 
    add: out std_logic_vector(3 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_50e644ef30;

architecture structural of add_convert1_entity_50e644ef30 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(3 downto 0);
  signal ce_1_sg_x338: std_logic;
  signal clk_1_sg_x338: std_logic;
  signal concat_y_net: std_logic_vector(4 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal delay13_q_net: std_logic_vector(3 downto 0);
  signal delay14_q_net: std_logic_vector(3 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(4 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(2 downto 0);
  signal new_add_y_net: std_logic_vector(3 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x338 <= ce_1;
  clk_1_sg_x338 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_8f12c32de0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 4,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 4,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x338,
      clk => clk_1_sg_x338,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_cf540617d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 5,
      y_width => 3
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 5,
      y_width => 4
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 5,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_42de9e04f9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(3 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_42de9e04f9;

architecture structural of cosin_entity_42de9e04f9 is
  signal assert_dout_net_x1: std_logic_vector(3 downto 0);
  signal ce_1_sg_x341: std_logic;
  signal clk_1_sg_x341: std_logic;
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(3 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x341 <= ce_1;
  clk_1_sg_x341 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_a9a42ddd37: entity work.add_convert0_entity_a9a42ddd37
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_50e644ef30: entity work.add_convert1_entity_50e644ef30
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 4,
      dout_width => 4
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x341,
      clk => clk_1_sg_x341,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x341,
      clk => clk_1_sg_x341,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x341,
      clk => clk_1_sg_x341,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_5e7b990fd3: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_467d752d46: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_core
    generic map (
      addr_width => 4,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_efdf1b1b05926829",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x341,
      a_clk => clk_1_sg_x341,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x341,
      b_clk => clk_1_sg_x341,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_8c5a8febd8 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_8c5a8febd8;

architecture structural of coeff_gen_entity_8c5a8febd8 is
  signal ce_1_sg_x342: std_logic;
  signal clk_1_sg_x342: std_logic;
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(3 downto 0);

begin
  ce_1_sg_x342 <= ce_1;
  clk_1_sg_x342 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_21d5d92029: entity work.bit_reverse_entity_21d5d92029
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_42de9e04f9: entity work.cosin_entity_42de9e04f9
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x342,
      clk => clk_1_sg_x342,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_f763d3ec59: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 11,
      x_width => 12,
      y_width => 4
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct/twiddle"

entity twiddle_entity_94bfa01a8b is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_94bfa01a8b;

architecture structural of twiddle_entity_94bfa01a8b is
  signal ce_1_sg_x343: std_logic;
  signal clk_1_sg_x343: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x343 <= ce_1;
  clk_1_sg_x343 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_a586ea121c: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x343,
      clk_1 => clk_1_sg_x343,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_9bfb22bcfc: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_bcb19b9074: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_926b2e72c1: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_099a550de5: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x343,
      clk_1 => clk_1_sg_x343,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_8c5a8febd8: entity work.coeff_gen_entity_8c5a8febd8
    port map (
      ce_1 => ce_1_sg_x343,
      clk_1 => clk_1_sg_x343,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/butterfly_direct"

entity butterfly_direct_entity_1af0b83f41 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_1af0b83f41;

architecture structural of butterfly_direct_entity_1af0b83f41 is
  signal ce_1_sg_x344: std_logic;
  signal clk_1_sg_x344: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x344 <= ce_1;
  clk_1_sg_x344 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_ff43c87dd4: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      dout => concatenate_y_net_x3
    );

  bus_convert_7be7051164: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_19dfb6c200: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_95b7493821: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_fbc223656a: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_67057968bb: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_f8c5fc3f6b: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_f9c2fe183f: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x344,
      clk => clk_1_sg_x344,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x344,
      clk => clk_1_sg_x344,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_9c8710f014: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x344,
      clk => clk_1_sg_x344,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_94bfa01a8b: entity work.twiddle_entity_94bfa01a8b
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x344,
      clk_1 => clk_1_sg_x344,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/delay_b"

entity delay_b_entity_00612e364c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_00612e364c;

architecture structural of delay_b_entity_00612e364c is
  signal ce_1_sg_x345: std_logic;
  signal clk_1_sg_x345: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x345 <= ce_1;
  clk_1_sg_x345 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 252,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_133a8817831fb97a",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x345,
      clk => clk_1_sg_x345,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 8,
      c_width => 36,
      core_name0 => "bmg_72_87bb354a843dab37",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x345,
      clk => clk_1_sg_x345,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5/sync_delay"

entity sync_delay_entity_a3a2369129 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_a3a2369129;

architecture structural of sync_delay_entity_a3a2369129 is
  signal ce_1_sg_x347: std_logic;
  signal clk_1_sg_x347: std_logic;
  signal constant1_op_net: std_logic_vector(8 downto 0);
  signal constant2_op_net: std_logic_vector(8 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(8 downto 0);
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x347 <= ce_1;
  clk_1_sg_x347 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_fd85eb7067
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_4a391b9a0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_b4ec9de7d1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_796a9d3dfbc0c498",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x347,
      clk => clk_1_sg_x347,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_6c3ee657fa
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_78eac2928d
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_5"

entity fft_stage_5_entity_14950a056d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_5_entity_14950a056d;

architecture structural of fft_stage_5_entity_14950a056d is
  signal ce_1_sg_x348: std_logic;
  signal clk_1_sg_x348: std_logic;
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x8: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x18: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x348 <= ce_1;
  clk_1_sg_x348 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x18 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x8 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x12;
  sync_out <= delay0_q_net_x3;

  butterfly_direct_1af0b83f41: entity work.butterfly_direct_entity_1af0b83f41
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x348,
      clk_1 => clk_1_sg_x348,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x12,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_12b8e0a4a9ef4845",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x348,
      clk => clk_1_sg_x348,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x2,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x348,
      clk => clk_1_sg_x348,
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => delay_q_net_x0
    );

  delay_b_00612e364c: entity work.delay_b_entity_00612e364c
    port map (
      ce_1 => ce_1_sg_x348,
      clk_1 => clk_1_sg_x348,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_a96c3f1545: entity work.delay_b_entity_00612e364c
    port map (
      ce_1 => ce_1_sg_x348,
      clk_1 => clk_1_sg_x348,
      din => reinterpret1_output_port_net_x18,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x348,
      clk => clk_1_sg_x348,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x348,
      clk => clk_1_sg_x348,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x3,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x348,
      clk => clk_1_sg_x348,
      clr => '0',
      d0 => reinterpret2_output_port_net_x3,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x8,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_a3a2369129: entity work.sync_delay_entity_a3a2369129
    port map (
      ce_1 => ce_1_sg_x348,
      clk_1 => clk_1_sg_x348,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_7c7c61e773 is
  port (
    in_x0: in std_logic_vector(4 downto 0); 
    out_x0: out std_logic_vector(4 downto 0)
  );
end bit_reverse_entity_7c7c61e773;

architecture structural of bit_reverse_entity_7c7c61e773 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(4 downto 0);
  signal slice_y_net_x0: std_logic_vector(4 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  concat: entity work.concat_2b3acb49f4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_3df356e0f9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(4 downto 0); 
    add: out std_logic_vector(4 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_3df356e0f9;

architecture structural of add_convert0_entity_3df356e0f9 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(4 downto 0);
  signal ce_1_sg_x375: std_logic;
  signal clk_1_sg_x375: std_logic;
  signal concat_y_net: std_logic_vector(5 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal delay13_q_net: std_logic_vector(4 downto 0);
  signal delay14_q_net: std_logic_vector(4 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(5 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(3 downto 0);
  signal new_add_y_net: std_logic_vector(4 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x375 <= ce_1;
  clk_1_sg_x375 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x375,
      clk => clk_1_sg_x375,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_ae3f02567e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 5,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 5,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x375,
      clk => clk_1_sg_x375,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x375,
      clk => clk_1_sg_x375,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x375,
      clk => clk_1_sg_x375,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x375,
      clk => clk_1_sg_x375,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_ac785d9b37
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 6,
      y_width => 4
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 6,
      y_width => 5
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 5,
      x_width => 6,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_a499587245 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(4 downto 0); 
    add: out std_logic_vector(4 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_a499587245;

architecture structural of add_convert1_entity_a499587245 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(4 downto 0);
  signal ce_1_sg_x376: std_logic;
  signal clk_1_sg_x376: std_logic;
  signal concat_y_net: std_logic_vector(5 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal delay13_q_net: std_logic_vector(4 downto 0);
  signal delay14_q_net: std_logic_vector(4 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(5 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(3 downto 0);
  signal new_add_y_net: std_logic_vector(4 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x376 <= ce_1;
  clk_1_sg_x376 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_ae3f02567e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 5,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 5,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x376,
      clk => clk_1_sg_x376,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_ac785d9b37
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 6,
      y_width => 4
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 6,
      y_width => 5
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 5,
      x_width => 6,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_299ac8b09e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(4 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_299ac8b09e;

architecture structural of cosin_entity_299ac8b09e is
  signal assert_dout_net_x1: std_logic_vector(4 downto 0);
  signal ce_1_sg_x379: std_logic;
  signal clk_1_sg_x379: std_logic;
  signal concat_y_net_x1: std_logic_vector(4 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(4 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x379 <= ce_1;
  clk_1_sg_x379 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_3df356e0f9: entity work.add_convert0_entity_3df356e0f9
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_a499587245: entity work.add_convert1_entity_a499587245
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 5,
      dout_width => 5
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x379,
      clk => clk_1_sg_x379,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x379,
      clk => clk_1_sg_x379,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x379,
      clk => clk_1_sg_x379,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_bd0d358d8c: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_3e07504796: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_core
    generic map (
      addr_width => 5,
      c_address_width => 5,
      c_width => 18,
      core_name0 => "dmg_72_1c323e86177437db",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x379,
      a_clk => clk_1_sg_x379,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x379,
      b_clk => clk_1_sg_x379,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_ba789e5070 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_ba789e5070;

architecture structural of coeff_gen_entity_ba789e5070 is
  signal ce_1_sg_x380: std_logic;
  signal clk_1_sg_x380: std_logic;
  signal concat_y_net_x1: std_logic_vector(4 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(4 downto 0);

begin
  ce_1_sg_x380 <= ce_1;
  clk_1_sg_x380 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_7c7c61e773: entity work.bit_reverse_entity_7c7c61e773
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_299ac8b09e: entity work.cosin_entity_299ac8b09e
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x380,
      clk => clk_1_sg_x380,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_cc8938b800: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 11,
      x_width => 12,
      y_width => 5
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct/twiddle"

entity twiddle_entity_07a2296890 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_07a2296890;

architecture structural of twiddle_entity_07a2296890 is
  signal ce_1_sg_x381: std_logic;
  signal clk_1_sg_x381: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x381 <= ce_1;
  clk_1_sg_x381 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_6a6baf78b5: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x381,
      clk_1 => clk_1_sg_x381,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_42db4e5a14: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_3ec198ae6d: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_5f87b43645: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_fe1bc13b0c: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x381,
      clk_1 => clk_1_sg_x381,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_ba789e5070: entity work.coeff_gen_entity_ba789e5070
    port map (
      ce_1 => ce_1_sg_x381,
      clk_1 => clk_1_sg_x381,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/butterfly_direct"

entity butterfly_direct_entity_d434e3f971 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_d434e3f971;

architecture structural of butterfly_direct_entity_d434e3f971 is
  signal ce_1_sg_x382: std_logic;
  signal clk_1_sg_x382: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x382 <= ce_1;
  clk_1_sg_x382 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_1360cc70be: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      dout => concatenate_y_net_x3
    );

  bus_convert_0b8dbfe466: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_f7b0c8beed: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_70945e41d2: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_01f541cdcb: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_4a0b12006b: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_667bd0db70: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_45df90e1ce: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x382,
      clk => clk_1_sg_x382,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x382,
      clk => clk_1_sg_x382,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_20ed3d3792: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x382,
      clk => clk_1_sg_x382,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_07a2296890: entity work.twiddle_entity_07a2296890
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x382,
      clk_1 => clk_1_sg_x382,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/delay_b"

entity delay_b_entity_497abae2ab is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_497abae2ab;

architecture structural of delay_b_entity_497abae2ab is
  signal ce_1_sg_x383: std_logic;
  signal clk_1_sg_x383: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x383 <= ce_1;
  clk_1_sg_x383 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 124,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_0c22adf9c6a5bc0d",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 7
    )
    port map (
      ce => ce_1_sg_x383,
      clk => clk_1_sg_x383,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 7,
      c_width => 36,
      core_name0 => "bmg_72_b92ee532c1b215f1",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x383,
      clk => clk_1_sg_x383,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6/sync_delay"

entity sync_delay_entity_85af25263b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_85af25263b;

architecture structural of sync_delay_entity_85af25263b is
  signal ce_1_sg_x385: std_logic;
  signal clk_1_sg_x385: std_logic;
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant2_op_net: std_logic_vector(7 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(7 downto 0);
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x385 <= ce_1;
  clk_1_sg_x385 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8aae5d3bb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_b437b02512
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_b7550dc611e0410a",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x385,
      clk => clk_1_sg_x385,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_54048c8b02
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_16235eb2bf
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_6"

entity fft_stage_6_entity_b55eecd3f6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_6_entity_b55eecd3f6;

architecture structural of fft_stage_6_entity_b55eecd3f6 is
  signal ce_1_sg_x386: std_logic;
  signal clk_1_sg_x386: std_logic;
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x9: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x386 <= ce_1;
  clk_1_sg_x386 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x14 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x9 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x15;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_d434e3f971: entity work.butterfly_direct_entity_d434e3f971
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x386,
      clk_1 => clk_1_sg_x386,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x15,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_133a8817831fb97a",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x386,
      clk => clk_1_sg_x386,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x4,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x386,
      clk => clk_1_sg_x386,
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => delay_q_net_x0
    );

  delay_b_497abae2ab: entity work.delay_b_entity_497abae2ab
    port map (
      ce_1 => ce_1_sg_x386,
      clk_1 => clk_1_sg_x386,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_1b5be235c4: entity work.delay_b_entity_497abae2ab
    port map (
      ce_1 => ce_1_sg_x386,
      clk_1 => clk_1_sg_x386,
      din => reinterpret1_output_port_net_x14,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x386,
      clk => clk_1_sg_x386,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x386,
      clk => clk_1_sg_x386,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x5,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x386,
      clk => clk_1_sg_x386,
      clr => '0',
      d0 => reinterpret2_output_port_net_x5,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x9,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_85af25263b: entity work.sync_delay_entity_85af25263b
    port map (
      ce_1 => ce_1_sg_x386,
      clk_1 => clk_1_sg_x386,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_d3a137e581 is
  port (
    in_x0: in std_logic_vector(5 downto 0); 
    out_x0: out std_logic_vector(5 downto 0)
  );
end bit_reverse_entity_d3a137e581;

architecture structural of bit_reverse_entity_d3a137e581 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(5 downto 0);
  signal slice_y_net_x0: std_logic_vector(5 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  concat: entity work.concat_2dc093ca7a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_d6ef9eb803 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(5 downto 0); 
    add: out std_logic_vector(5 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_d6ef9eb803;

architecture structural of add_convert0_entity_d6ef9eb803 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(5 downto 0);
  signal ce_1_sg_x413: std_logic;
  signal clk_1_sg_x413: std_logic;
  signal concat_y_net: std_logic_vector(6 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(5 downto 0);
  signal delay13_q_net: std_logic_vector(5 downto 0);
  signal delay14_q_net: std_logic_vector(5 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(6 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(4 downto 0);
  signal new_add_y_net: std_logic_vector(5 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x413 <= ce_1;
  clk_1_sg_x413 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x413,
      clk => clk_1_sg_x413,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_75261c7c53
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 6,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 6,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x413,
      clk => clk_1_sg_x413,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_0b18d34058
    port map (
      ce => ce_1_sg_x413,
      clk => clk_1_sg_x413,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_0b18d34058
    port map (
      ce => ce_1_sg_x413,
      clk => clk_1_sg_x413,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x413,
      clk => clk_1_sg_x413,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 7,
      y_width => 5
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 7,
      y_width => 6
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 7,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_96d1ac614c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(5 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_96d1ac614c;

architecture structural of add_convert1_entity_96d1ac614c is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(5 downto 0);
  signal ce_1_sg_x414: std_logic;
  signal clk_1_sg_x414: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(6 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x414 <= ce_1;
  clk_1_sg_x414 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x414,
      clk => clk_1_sg_x414,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x414,
      clk => clk_1_sg_x414,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x414,
      clk => clk_1_sg_x414,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 7,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_5c7a19b8b5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(5 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_5c7a19b8b5;

architecture structural of cosin_entity_5c7a19b8b5 is
  signal assert_dout_net_x1: std_logic_vector(5 downto 0);
  signal ce_1_sg_x417: std_logic;
  signal clk_1_sg_x417: std_logic;
  signal concat_y_net_x1: std_logic_vector(5 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(5 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x417 <= ce_1;
  clk_1_sg_x417 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_d6ef9eb803: entity work.add_convert0_entity_d6ef9eb803
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_96d1ac614c: entity work.add_convert1_entity_96d1ac614c
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 6,
      dout_width => 6
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_d976c6caad: entity work.c_to_ri_entity_8f95d0368d
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x417,
      clk => clk_1_sg_x417,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x417,
      clk => clk_1_sg_x417,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x417,
      clk => clk_1_sg_x417,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_f5f95aec2d: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_69d8c6c193: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_core
    generic map (
      c_address_width => 6,
      c_width => 36,
      core_name0 => "bmg_72_eb304381eda4ae1e",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x417,
      clk => clk_1_sg_x417,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_ba6ec8207d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_ba6ec8207d;

architecture structural of coeff_gen_entity_ba6ec8207d is
  signal ce_1_sg_x418: std_logic;
  signal clk_1_sg_x418: std_logic;
  signal concat_y_net_x1: std_logic_vector(5 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x418 <= ce_1;
  clk_1_sg_x418 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_d3a137e581: entity work.bit_reverse_entity_d3a137e581
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_5c7a19b8b5: entity work.cosin_entity_5c7a19b8b5
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x418,
      clk => clk_1_sg_x418,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_ca5672875d: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 11,
      x_width => 12,
      y_width => 6
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct/twiddle"

entity twiddle_entity_1cb59b1c90 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_1cb59b1c90;

architecture structural of twiddle_entity_1cb59b1c90 is
  signal ce_1_sg_x419: std_logic;
  signal clk_1_sg_x419: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x419 <= ce_1;
  clk_1_sg_x419 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_416dbe56c8: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x419,
      clk_1 => clk_1_sg_x419,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_4c0748d19f: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_2e688f71a3: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_fc01e4026c: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_eeb4398156: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x419,
      clk_1 => clk_1_sg_x419,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_ba6ec8207d: entity work.coeff_gen_entity_ba6ec8207d
    port map (
      ce_1 => ce_1_sg_x419,
      clk_1 => clk_1_sg_x419,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/butterfly_direct"

entity butterfly_direct_entity_48daf0a77b is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_48daf0a77b;

architecture structural of butterfly_direct_entity_48daf0a77b is
  signal ce_1_sg_x420: std_logic;
  signal clk_1_sg_x420: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x420 <= ce_1;
  clk_1_sg_x420 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_b6ec5dd49a: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      dout => concatenate_y_net_x3
    );

  bus_convert_bc8eab82b7: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_92496074de: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_200d65fc8f: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_c8af661677: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_1a0fb95990: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_c62f398c73: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_e1678a56ee: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x420,
      clk => clk_1_sg_x420,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x420,
      clk => clk_1_sg_x420,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_63f70a4285: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x420,
      clk => clk_1_sg_x420,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_1cb59b1c90: entity work.twiddle_entity_1cb59b1c90
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x420,
      clk_1 => clk_1_sg_x420,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/delay_b"

entity delay_b_entity_55888c2f28 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_55888c2f28;

architecture structural of delay_b_entity_55888c2f28 is
  signal ce_1_sg_x421: std_logic;
  signal clk_1_sg_x421: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x421 <= ce_1;
  clk_1_sg_x421 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 60,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_d60ecc44fc05ecdd",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x421,
      clk => clk_1_sg_x421,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 6,
      c_width => 36,
      core_name0 => "bmg_72_59143b4ed22b761d",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x421,
      clk => clk_1_sg_x421,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7/sync_delay"

entity sync_delay_entity_fec4c0d8d2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_fec4c0d8d2;

architecture structural of sync_delay_entity_fec4c0d8d2 is
  signal ce_1_sg_x423: std_logic;
  signal clk_1_sg_x423: std_logic;
  signal constant1_op_net: std_logic_vector(6 downto 0);
  signal constant2_op_net: std_logic_vector(6 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(6 downto 0);
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x423 <= ce_1;
  clk_1_sg_x423 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_7244cd602b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_7b07120b87
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_180df391de
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_03f06ae367a98e8a",
      op_arith => xlUnsigned,
      op_width => 7
    )
    port map (
      ce => ce_1_sg_x423,
      clk => clk_1_sg_x423,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_9a3978c602
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_23065a6aa3
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_7"

entity fft_stage_7_entity_c4300ce589 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_7_entity_c4300ce589;

architecture structural of fft_stage_7_entity_c4300ce589 is
  signal ce_1_sg_x424: std_logic;
  signal clk_1_sg_x424: std_logic;
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x10: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x424 <= ce_1;
  clk_1_sg_x424 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x17 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x10 <= shift;
  delay0_q_net_x6 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x12;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_48daf0a77b: entity work.butterfly_direct_entity_48daf0a77b
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x424,
      clk_1 => clk_1_sg_x424,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x12,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_0c22adf9c6a5bc0d",
      op_arith => xlUnsigned,
      op_width => 7
    )
    port map (
      ce => ce_1_sg_x424,
      clk => clk_1_sg_x424,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x6,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x424,
      clk => clk_1_sg_x424,
      clr => '0',
      d(0) => delay0_q_net_x6,
      q(0) => delay_q_net_x0
    );

  delay_b_55888c2f28: entity work.delay_b_entity_55888c2f28
    port map (
      ce_1 => ce_1_sg_x424,
      clk_1 => clk_1_sg_x424,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_4e132ccc01: entity work.delay_b_entity_55888c2f28
    port map (
      ce_1 => ce_1_sg_x424,
      clk_1 => clk_1_sg_x424,
      din => reinterpret1_output_port_net_x17,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x424,
      clk => clk_1_sg_x424,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x424,
      clk => clk_1_sg_x424,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x7,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x424,
      clk => clk_1_sg_x424,
      clr => '0',
      d0 => reinterpret2_output_port_net_x7,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x10,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_fec4c0d8d2: entity work.sync_delay_entity_fec4c0d8d2
    port map (
      ce_1 => ce_1_sg_x424,
      clk_1 => clk_1_sg_x424,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_abec178d91 is
  port (
    in_x0: in std_logic_vector(6 downto 0); 
    out_x0: out std_logic_vector(6 downto 0)
  );
end bit_reverse_entity_abec178d91;

architecture structural of bit_reverse_entity_abec178d91 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(6 downto 0);
  signal slice_y_net_x0: std_logic_vector(6 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  concat: entity work.concat_eb5f1ca7f9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_f1edfbee00 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(6 downto 0); 
    add: out std_logic_vector(6 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_f1edfbee00;

architecture structural of add_convert0_entity_f1edfbee00 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(6 downto 0);
  signal ce_1_sg_x451: std_logic;
  signal clk_1_sg_x451: std_logic;
  signal concat_y_net: std_logic_vector(7 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(6 downto 0);
  signal delay13_q_net: std_logic_vector(6 downto 0);
  signal delay14_q_net: std_logic_vector(6 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(7 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(5 downto 0);
  signal new_add_y_net: std_logic_vector(6 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x451 <= ce_1;
  clk_1_sg_x451 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x451,
      clk => clk_1_sg_x451,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_dc245eb1d2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 7,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 7,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x451,
      clk => clk_1_sg_x451,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_9066adfc41
    port map (
      ce => ce_1_sg_x451,
      clk => clk_1_sg_x451,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_9066adfc41
    port map (
      ce => ce_1_sg_x451,
      clk => clk_1_sg_x451,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x451,
      clk => clk_1_sg_x451,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_83e473517e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 6,
      x_width => 8,
      y_width => 7
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 7,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_7c29727ce3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(6 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_7c29727ce3;

architecture structural of add_convert1_entity_7c29727ce3 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(6 downto 0);
  signal ce_1_sg_x452: std_logic;
  signal clk_1_sg_x452: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(7 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x452 <= ce_1;
  clk_1_sg_x452 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x452,
      clk => clk_1_sg_x452,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x452,
      clk => clk_1_sg_x452,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x452,
      clk => clk_1_sg_x452,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_83e473517e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 7,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_36999f42d0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(6 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_36999f42d0;

architecture structural of cosin_entity_36999f42d0 is
  signal assert_dout_net_x1: std_logic_vector(6 downto 0);
  signal ce_1_sg_x455: std_logic;
  signal clk_1_sg_x455: std_logic;
  signal concat_y_net_x1: std_logic_vector(6 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(6 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x455 <= ce_1;
  clk_1_sg_x455 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_f1edfbee00: entity work.add_convert0_entity_f1edfbee00
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_7c29727ce3: entity work.add_convert1_entity_7c29727ce3
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 7,
      dout_width => 7
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_82f5294717: entity work.c_to_ri_entity_8f95d0368d
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x455,
      clk => clk_1_sg_x455,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x455,
      clk => clk_1_sg_x455,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x455,
      clk => clk_1_sg_x455,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_cc3fc2206a: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_4b8f331d6e: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_core
    generic map (
      c_address_width => 7,
      c_width => 36,
      core_name0 => "bmg_72_6711bf92f3a48934",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x455,
      clk => clk_1_sg_x455,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_981aec6c3a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_981aec6c3a;

architecture structural of coeff_gen_entity_981aec6c3a is
  signal ce_1_sg_x456: std_logic;
  signal clk_1_sg_x456: std_logic;
  signal concat_y_net_x1: std_logic_vector(6 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(6 downto 0);

begin
  ce_1_sg_x456 <= ce_1;
  clk_1_sg_x456 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_abec178d91: entity work.bit_reverse_entity_abec178d91
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_36999f42d0: entity work.cosin_entity_36999f42d0
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x456,
      clk => clk_1_sg_x456,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_3a7e601112: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 11,
      x_width => 12,
      y_width => 7
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct/twiddle"

entity twiddle_entity_d9466e5aba is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_d9466e5aba;

architecture structural of twiddle_entity_d9466e5aba is
  signal ce_1_sg_x457: std_logic;
  signal clk_1_sg_x457: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal ram_data_out_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  ram_data_out_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x457 <= ce_1;
  clk_1_sg_x457 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_0651c23458: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x457,
      clk_1 => clk_1_sg_x457,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_c860c7035c: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => ram_data_out_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_c0d50050c9: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_ec93fef2c7: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_81dd5502ad: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x457,
      clk_1 => clk_1_sg_x457,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_981aec6c3a: entity work.coeff_gen_entity_981aec6c3a
    port map (
      ce_1 => ce_1_sg_x457,
      clk_1 => clk_1_sg_x457,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/butterfly_direct"

entity butterfly_direct_entity_be50e176da is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_be50e176da;

architecture structural of butterfly_direct_entity_be50e176da is
  signal ce_1_sg_x458: std_logic;
  signal clk_1_sg_x458: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay2_q_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ram_data_out_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x458 <= ce_1;
  clk_1_sg_x458 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x0;

  bus_add_1674bd58c4: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      dout => concatenate_y_net_x3
    );

  bus_convert_b31030a14b: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_6d91e9f1c1: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_12c2dd663d: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_46c6eb5557: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_12e44be69b: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_b5532f9ecf: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_1aca6c843c: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x458,
      clk => clk_1_sg_x458,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x458,
      clk => clk_1_sg_x458,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_5b68c973fe: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x458,
      clk => clk_1_sg_x458,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_d9466e5aba: entity work.twiddle_entity_d9466e5aba
    port map (
      ai => ram_data_out_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x458,
      clk_1 => clk_1_sg_x458,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/delay_b"

entity delay_b_entity_4bce676126 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_4bce676126;

architecture structural of delay_b_entity_4bce676126 is
  signal ce_1_sg_x459: std_logic;
  signal clk_1_sg_x459: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(4 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x459 <= ce_1;
  clk_1_sg_x459 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= ram_data_out_net_x3;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.xlcounter_limit_fft_core
    generic map (
      cnt_15_0 => 28,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_ee60311bb9d0db53",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 5
    )
    port map (
      ce => ce_1_sg_x459,
      clk => clk_1_sg_x459,
      clr => '0',
      en => "1",
      rst => "0",
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_core
    generic map (
      c_address_width => 5,
      c_width => 36,
      core_name0 => "bmg_72_ba1afd1a3b6d9138",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x459,
      clk => clk_1_sg_x459,
      data_in => mux1_y_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8/sync_delay"

entity sync_delay_entity_ee87732189 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_ee87732189;

architecture structural of sync_delay_entity_ee87732189 is
  signal ce_1_sg_x461: std_logic;
  signal clk_1_sg_x461: std_logic;
  signal constant1_op_net: std_logic_vector(5 downto 0);
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(5 downto 0);
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x461 <= ce_1;
  clk_1_sg_x461 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_7ea0f2fff7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_961b61f8a1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a267c870be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_cb1ffe90ceffe54f",
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x461,
      clk => clk_1_sg_x461,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_931d61fb72
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_fe487ce1c7
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_8"

entity fft_stage_8_entity_518409c227 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_8_entity_518409c227;

architecture structural of fft_stage_8_entity_518409c227 is
  signal ce_1_sg_x462: std_logic;
  signal clk_1_sg_x462: std_logic;
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fft_shift_net_x11: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x462 <= ce_1;
  clk_1_sg_x462 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x14 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x11 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x15;
  sync_out <= delay0_q_net_x3;

  butterfly_direct_be50e176da: entity work.butterfly_direct_entity_be50e176da
    port map (
      a => ram_data_out_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x462,
      clk_1 => clk_1_sg_x462,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x15,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_d60ecc44fc05ecdd",
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x462,
      clk => clk_1_sg_x462,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x2,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x462,
      clk => clk_1_sg_x462,
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => delay_q_net_x0
    );

  delay_b_4bce676126: entity work.delay_b_entity_4bce676126
    port map (
      ce_1 => ce_1_sg_x462,
      clk_1 => clk_1_sg_x462,
      din => mux1_y_net_x0,
      dout => ram_data_out_net_x3
    );

  delay_f_87a6813b24: entity work.delay_b_entity_4bce676126
    port map (
      ce_1 => ce_1_sg_x462,
      clk_1 => clk_1_sg_x462,
      din => reinterpret1_output_port_net_x14,
      dout => ram_data_out_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x462,
      clk => clk_1_sg_x462,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x462,
      clk => clk_1_sg_x462,
      clr => '0',
      d0 => ram_data_out_net_x0,
      d1 => reinterpret2_output_port_net_x3,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x462,
      clk => clk_1_sg_x462,
      clr => '0',
      d0 => reinterpret2_output_port_net_x3,
      d1 => ram_data_out_net_x0,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x11,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_ee87732189: entity work.sync_delay_entity_ee87732189
    port map (
      ce_1 => ce_1_sg_x462,
      clk_1 => clk_1_sg_x462,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_e98cf63321 is
  port (
    in_x0: in std_logic_vector(7 downto 0); 
    out_x0: out std_logic_vector(7 downto 0)
  );
end bit_reverse_entity_e98cf63321;

architecture structural of bit_reverse_entity_e98cf63321 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal slice_y_net_x0: std_logic_vector(7 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  concat: entity work.concat_7673b9b993
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_8f9be6a1fa is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(7 downto 0); 
    add: out std_logic_vector(7 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_8f9be6a1fa;

architecture structural of add_convert0_entity_8f9be6a1fa is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(7 downto 0);
  signal ce_1_sg_x489: std_logic;
  signal clk_1_sg_x489: std_logic;
  signal concat_y_net: std_logic_vector(8 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(7 downto 0);
  signal delay13_q_net: std_logic_vector(7 downto 0);
  signal delay14_q_net: std_logic_vector(7 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(8 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(6 downto 0);
  signal new_add_y_net: std_logic_vector(7 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x489 <= ce_1;
  clk_1_sg_x489 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x489,
      clk => clk_1_sg_x489,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  concat: entity work.concat_f62149b02a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 8,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 8,
      latency => 1,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x489,
      clk => clk_1_sg_x489,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_ebec135d8a
    port map (
      ce => ce_1_sg_x489,
      clk => clk_1_sg_x489,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_ebec135d8a
    port map (
      ce => ce_1_sg_x489,
      clk => clk_1_sg_x489,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x489,
      clk => clk_1_sg_x489,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_1ece14600f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 6,
      x_width => 9,
      y_width => 7
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 9,
      y_width => 8
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 8,
      x_width => 9,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_870a0a1d4c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(7 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_870a0a1d4c;

architecture structural of add_convert1_entity_870a0a1d4c is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x490: std_logic;
  signal clk_1_sg_x490: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(8 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x490 <= ce_1;
  clk_1_sg_x490 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.xladdsub_fft_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 2,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 2,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 3,
      core_name0 => "addsb_11_0_c8fdf7c1ceafa9d8",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 3,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 2
    )
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x490,
      clk => clk_1_sg_x490,
      clr => '0',
      en => "1",
      s => addsub5_s_net
    );

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x490,
      clk => clk_1_sg_x490,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x490,
      clk => clk_1_sg_x490,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_1ece14600f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 8,
      x_width => 9,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_7a3faf875c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(7 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_7a3faf875c;

architecture structural of cosin_entity_7a3faf875c is
  signal assert_dout_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x493: std_logic;
  signal clk_1_sg_x493: std_logic;
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(7 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x493 <= ce_1;
  clk_1_sg_x493 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_8f9be6a1fa: entity work.add_convert0_entity_8f9be6a1fa
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_870a0a1d4c: entity work.add_convert1_entity_870a0a1d4c
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 8,
      dout_width => 8
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_b4455b1101: entity work.c_to_ri_entity_8f95d0368d
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x493,
      clk => clk_1_sg_x493,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x493,
      clk => clk_1_sg_x493,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x493,
      clk => clk_1_sg_x493,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_ce7898510f: entity work.invert0_entity_e94ce56a25
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_302423a94b: entity work.invert1_entity_56100eb48e
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_core
    generic map (
      c_address_width => 8,
      c_width => 36,
      core_name0 => "bmg_72_070de696ab472038",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x493,
      clk => clk_1_sg_x493,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_e5446135f7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_e5446135f7;

architecture structural of coeff_gen_entity_e5446135f7 is
  signal ce_1_sg_x494: std_logic;
  signal clk_1_sg_x494: std_logic;
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal mux_y_net_x6: std_logic;
  signal slice_y_net_x0: std_logic_vector(7 downto 0);

begin
  ce_1_sg_x494 <= ce_1;
  clk_1_sg_x494 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x6 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_e98cf63321: entity work.bit_reverse_entity_e98cf63321
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_7a3faf875c: entity work.cosin_entity_7a3faf875c
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ed810b6704650710",
      op_arith => xlUnsigned,
      op_width => 12
    )
    port map (
      ce => ce_1_sg_x494,
      clk => clk_1_sg_x494,
      clr => '0',
      en => "1",
      rst(0) => mux_y_net_x6,
      op => counter_op_net
    );

  ri_to_c_3b14128470: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 11,
      x_width => 12,
      y_width => 8
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct/twiddle"

entity twiddle_entity_37a13b45f1 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_37a13b45f1;

architecture structural of twiddle_entity_37a13b45f1 is
  signal ce_1_sg_x495: std_logic;
  signal clk_1_sg_x495: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal delay_q_net_x1: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal mux_y_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x7: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  delay_q_net_x1 <= ai;
  mux_y_net_x2 <= bi;
  ce_1_sg_x495 <= ce_1;
  clk_1_sg_x495 <= clk_1;
  mux_y_net_x7 <= sync_in;
  ao <= reinterpret1_output_port_net_x10;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_77e2c1cf91: entity work.bus_convert_entity_a82e0e1650
    port map (
      ce_1 => ce_1_sg_x495,
      clk_1 => clk_1_sg_x495,
      din => reinterpret1_output_port_net_x9,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_54042430b5: entity work.bus_create_entity_9c2c0dccf0
    port map (
      in1 => mux_y_net_x2,
      in2 => mux_y_net_x7,
      in3 => delay_q_net_x1,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_97d349be3c: entity work.bus_expand1_entity_e394667c48
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x10,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_80272b418b: entity work.bus_expand_entity_ad772b3d60
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x8,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_c982f7443c: entity work.bus_mult_entity_f9d9d4b2f7
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x495,
      clk_1 => clk_1_sg_x495,
      misci => reinterpret1_output_port_net_x8,
      a_b => reinterpret1_output_port_net_x9,
      misco => dmisc_q_net_x2
    );

  coeff_gen_e5446135f7: entity work.coeff_gen_entity_e5446135f7
    port map (
      ce_1 => ce_1_sg_x495,
      clk_1 => clk_1_sg_x495,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x7,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/butterfly_direct"

entity butterfly_direct_entity_df7b28d60f is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_df7b28d60f;

architecture structural of butterfly_direct_entity_df7b28d60f is
  signal ce_1_sg_x496: std_logic;
  signal clk_1_sg_x496: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay2_q_net: std_logic;
  signal delay_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic_vector(83 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x8: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice2_y_net_x1: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  delay_q_net_x2 <= a;
  mux_y_net_x3 <= b;
  ce_1_sg_x496 <= ce_1;
  clk_1_sg_x496 <= clk_1;
  slice_y_net_x0 <= shift;
  mux_y_net_x8 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x2;
  of_x0 <= reinterpret1_output_port_net_x11;
  sync_out <= delay0_q_net_x2;

  bus_add_ed66ecf2db: entity work.bus_add_entity_fda2dbc1e4
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      dout => concatenate_y_net_x3
    );

  bus_convert_d8feef432d: entity work.bus_convert_entity_b21c3d5983
    port map (
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      din => mux_y_net_x1,
      dout => concatenate_y_net_x4,
      overflow => concatenate_y_net_x5
    );

  bus_expand_cb96dd5627: entity work.bus_expand_entity_2ff4545d65
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x2
    );

  bus_norm0_b2807d9fab: entity work.bus_norm0_entity_19ac017aaf
    port map (
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x1
    );

  bus_norm1_15baeee458: entity work.bus_norm1_entity_d801aceba7
    port map (
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      din => concatenate_y_net_x7,
      dout => concatenate_y_net_x6
    );

  bus_relational_59772c7020: entity work.bus_relational_entity_53f1d0be84
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x11
    );

  bus_scale_0d602ef32b: entity work.bus_scale_entity_cc780061b4
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_sub_d41b2631cb: entity work.bus_sub_entity_5f1ccce5f7
    port map (
      a => reinterpret1_output_port_net_x10,
      b => concatenate_y_net_x9,
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      dout => concatenate_y_net_x8
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x8,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x496,
      clk => clk_1_sg_x496,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x2
    );

  delay2: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x496,
      clk => clk_1_sg_x496,
      clr => '0',
      d(0) => slice_y_net_x0,
      q(0) => delay2_q_net
    );

  munge_f7ee95b389: entity work.munge_entity_597456506f
    port map (
      din => concatenate_y_net_x5,
      dout => reinterpret_out_output_port_net_x2
    );

  mux: entity work.mux_86d5838e9c
    port map (
      ce => ce_1_sg_x496,
      clk => clk_1_sg_x496,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => concatenate_y_net_x6,
      sel(0) => delay2_q_net,
      y => mux_y_net_x1
    );

  twiddle_37a13b45f1: entity work.twiddle_entity_37a13b45f1
    port map (
      ai => delay_q_net_x2,
      bi => mux_y_net_x3,
      ce_1 => ce_1_sg_x496,
      clk_1 => clk_1_sg_x496,
      sync_in => mux_y_net_x8,
      ao => reinterpret1_output_port_net_x10,
      bwo => concatenate_y_net_x9,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/delay_b"

entity delay_b_entity_8d0a68a4c7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay_b_entity_8d0a68a4c7;

architecture structural of delay_b_entity_8d0a68a4c7 is
  signal ce_1_sg_x497: std_logic;
  signal clk_1_sg_x497: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x497 <= ce_1;
  clk_1_sg_x497 <= clk_1;
  mux1_y_net_x0 <= din;
  dout <= delay_q_net_x3;

  delay: entity work.delay_3a3620b5a6
    port map (
      ce => ce_1_sg_x497,
      clk => clk_1_sg_x497,
      clr => '0',
      d => mux1_y_net_x0,
      q => delay_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9/sync_delay"

entity sync_delay_entity_605dfe71ca is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_605dfe71ca;

architecture structural of sync_delay_entity_605dfe71ca is
  signal ce_1_sg_x499: std_logic;
  signal clk_1_sg_x499: std_logic;
  signal constant1_op_net: std_logic_vector(4 downto 0);
  signal constant2_op_net: std_logic_vector(4 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(4 downto 0);
  signal counter_op_net: std_logic_vector(4 downto 0);
  signal delay_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x9: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x499 <= ce_1;
  clk_1_sg_x499 <= clk_1;
  delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x9;

  constant1: entity work.constant_fe72737ca0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_ef0e2e5fc6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_582a3706dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_d5eedfa744d4da30",
      op_arith => xlUnsigned,
      op_width => 5
    )
    port map (
      ce => ce_1_sg_x499,
      clk => clk_1_sg_x499,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => delay_q_net_x0,
      rst => "0",
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x9
    );

  relational: entity work.relational_9ece3c8c4e
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_dc5bc996c9
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core/fft_stage_9"

entity fft_stage_9_entity_f8166671d4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_9_entity_f8166671d4;

architecture structural of fft_stage_9_entity_f8166671d4 is
  signal ce_1_sg_x500: std_logic;
  signal clk_1_sg_x500: std_logic;
  signal counter_op_net: std_logic_vector(4 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay_q_net_x0: std_logic;
  signal delay_q_net_x3: std_logic_vector(35 downto 0);
  signal delay_q_net_x4: std_logic_vector(35 downto 0);
  signal fft_shift_net_x12: std_logic_vector(31 downto 0);
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic_vector(35 downto 0);
  signal mux_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice_y_net_x0: std_logic;

begin
  ce_1_sg_x500 <= ce_1;
  clk_1_sg_x500 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x17 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x12 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x4;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x12;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_df7b28d60f: entity work.butterfly_direct_entity_df7b28d60f
    port map (
      a => delay_q_net_x3,
      b => mux_y_net_x3,
      ce_1 => ce_1_sg_x500,
      clk_1 => clk_1_sg_x500,
      shift => slice_y_net_x0,
      sync_in => mux_y_net_x9,
      a_bw => reinterpret1_output_port_net_x12,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.xlcounter_free_fft_core
    generic map (
      core_name0 => "cntr_11_0_ee60311bb9d0db53",
      op_arith => xlUnsigned,
      op_width => 5
    )
    port map (
      ce => ce_1_sg_x500,
      clk => clk_1_sg_x500,
      clr => '0',
      en => "1",
      rst(0) => delay0_q_net_x4,
      op => counter_op_net
    );

  delay: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x500,
      clk => clk_1_sg_x500,
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => delay_q_net_x0
    );

  delay_b_8d0a68a4c7: entity work.delay_b_entity_8d0a68a4c7
    port map (
      ce_1 => ce_1_sg_x500,
      clk_1 => clk_1_sg_x500,
      din => mux1_y_net_x0,
      dout => delay_q_net_x3
    );

  delay_f_9a5d319ac1: entity work.delay_b_entity_8d0a68a4c7
    port map (
      ce_1 => ce_1_sg_x500,
      clk_1 => clk_1_sg_x500,
      din => reinterpret1_output_port_net_x17,
      dout => delay_q_net_x4
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x500,
      clk => clk_1_sg_x500,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x11,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x4
    );

  mux: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x500,
      clk => clk_1_sg_x500,
      clr => '0',
      d0 => delay_q_net_x4,
      d1 => reinterpret2_output_port_net_x5,
      sel(0) => slice1_y_net,
      y => mux_y_net_x3
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x500,
      clk => clk_1_sg_x500,
      clr => '0',
      d0 => reinterpret2_output_port_net_x5,
      d1 => delay_q_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x12,
      y(0) => slice_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_605dfe71ca: entity work.sync_delay_entity_605dfe71ca
    port map (
      ce_1 => ce_1_sg_x500,
      clk_1 => clk_1_sg_x500,
      in_x0 => delay_q_net_x0,
      out_x0 => mux_y_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2/biplex_core"

entity biplex_core_entity_a39782552e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    pol1: in std_logic_vector(35 downto 0); 
    pol2: in std_logic_vector(35 downto 0); 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end biplex_core_entity_a39782552e;

architecture structural of biplex_core_entity_a39782552e is
  signal ce_1_sg_x501: std_logic;
  signal clk_1_sg_x501: std_logic;
  signal constant_op_net_x0: std_logic;
  signal delay0_q_net_x10: std_logic;
  signal delay0_q_net_x11: std_logic;
  signal delay0_q_net_x12: std_logic;
  signal delay0_q_net_x13: std_logic;
  signal delay0_q_net_x14: std_logic;
  signal delay0_q_net_x15: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal delay0_q_net_x7: std_logic;
  signal delay0_q_net_x8: std_logic;
  signal delay0_q_net_x9: std_logic;
  signal fft_shift_net_x13: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x10: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x12: std_logic;
  signal logical1_y_net_x13: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical1_y_net_x7: std_logic;
  signal logical1_y_net_x8: std_logic;
  signal logical1_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x18: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x19: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x20: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x21: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x22: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x23: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x24: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x25: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x26: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x27: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x13: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x9: std_logic_vector(35 downto 0);
  signal sync_net_x1: std_logic;

begin
  ce_1_sg_x501 <= ce_1;
  clk_1_sg_x501 <= clk_1;
  reinterpret1_output_port_net_x16 <= pol1;
  reinterpret1_output_port_net_x26 <= pol2;
  fft_shift_net_x13 <= shift;
  sync_net_x1 <= sync;
  of_x0 <= logical1_y_net_x13;
  out1 <= reinterpret2_output_port_net_x16;
  out2 <= reinterpret1_output_port_net_x27;
  sync_out <= delay0_q_net_x15;

  constant_x0: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net_x0
    );

  fft_stage_10_3b39e0a900: entity work.fft_stage_10_entity_3b39e0a900
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x6,
      in2 => reinterpret1_output_port_net_x25,
      of_in => logical1_y_net_x12,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x14,
      of_x0 => logical1_y_net_x3,
      out1 => reinterpret2_output_port_net_x4,
      out2 => reinterpret1_output_port_net_x14,
      sync_out => delay0_q_net_x3
    );

  fft_stage_11_4f6b9006ee: entity work.fft_stage_11_entity_4f6b9006ee
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x4,
      in2 => reinterpret1_output_port_net_x14,
      of_in => logical1_y_net_x3,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x3,
      of_x0 => logical1_y_net_x2,
      out1 => reinterpret2_output_port_net_x5,
      out2 => reinterpret1_output_port_net_x17,
      sync_out => delay0_q_net_x5
    );

  fft_stage_12_4d66daf6cf: entity work.fft_stage_12_entity_4d66daf6cf
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x5,
      in2 => reinterpret1_output_port_net_x17,
      of_in => logical1_y_net_x2,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x5,
      of_x0 => logical1_y_net_x4,
      out1 => reinterpret2_output_port_net_x7,
      out2 => reinterpret1_output_port_net_x18,
      sync_out => delay0_q_net_x6
    );

  fft_stage_13_02afd91842: entity work.fft_stage_13_entity_02afd91842
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x7,
      in2 => reinterpret1_output_port_net_x18,
      of_in => logical1_y_net_x4,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x6,
      of_x0 => logical1_y_net_x13,
      out1 => reinterpret2_output_port_net_x16,
      out2 => reinterpret1_output_port_net_x27,
      sync_out => delay0_q_net_x15
    );

  fft_stage_1_a0aa893753: entity work.fft_stage_1_entity_a0aa893753
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret1_output_port_net_x16,
      in2 => reinterpret1_output_port_net_x26,
      of_in => constant_op_net_x0,
      shift => fft_shift_net_x13,
      sync => sync_net_x1,
      of_x0 => logical1_y_net_x1,
      out1 => reinterpret2_output_port_net_x3,
      out2 => reinterpret1_output_port_net_x8,
      sync_out => delay0_q_net_x2
    );

  fft_stage_2_012e00c14b: entity work.fft_stage_2_entity_012e00c14b
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x3,
      in2 => reinterpret1_output_port_net_x8,
      of_in => logical1_y_net_x1,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x2,
      of_x0 => logical1_y_net_x5,
      out1 => reinterpret2_output_port_net_x9,
      out2 => reinterpret1_output_port_net_x12,
      sync_out => delay0_q_net_x7
    );

  fft_stage_3_33ea5e4989: entity work.fft_stage_3_entity_33ea5e4989
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x9,
      in2 => reinterpret1_output_port_net_x12,
      of_in => logical1_y_net_x5,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x7,
      of_x0 => logical1_y_net_x6,
      out1 => reinterpret2_output_port_net_x10,
      out2 => reinterpret1_output_port_net_x19,
      sync_out => delay0_q_net_x8
    );

  fft_stage_4_a779b0edc3: entity work.fft_stage_4_entity_a779b0edc3
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x10,
      in2 => reinterpret1_output_port_net_x19,
      of_in => logical1_y_net_x6,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x8,
      of_x0 => logical1_y_net_x7,
      out1 => reinterpret2_output_port_net_x11,
      out2 => reinterpret1_output_port_net_x20,
      sync_out => delay0_q_net_x9
    );

  fft_stage_5_14950a056d: entity work.fft_stage_5_entity_14950a056d
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x11,
      in2 => reinterpret1_output_port_net_x20,
      of_in => logical1_y_net_x7,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x9,
      of_x0 => logical1_y_net_x8,
      out1 => reinterpret2_output_port_net_x12,
      out2 => reinterpret1_output_port_net_x21,
      sync_out => delay0_q_net_x10
    );

  fft_stage_6_b55eecd3f6: entity work.fft_stage_6_entity_b55eecd3f6
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x12,
      in2 => reinterpret1_output_port_net_x21,
      of_in => logical1_y_net_x8,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x10,
      of_x0 => logical1_y_net_x9,
      out1 => reinterpret2_output_port_net_x13,
      out2 => reinterpret1_output_port_net_x22,
      sync_out => delay0_q_net_x11
    );

  fft_stage_7_c4300ce589: entity work.fft_stage_7_entity_c4300ce589
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x13,
      in2 => reinterpret1_output_port_net_x22,
      of_in => logical1_y_net_x9,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x11,
      of_x0 => logical1_y_net_x10,
      out1 => reinterpret2_output_port_net_x14,
      out2 => reinterpret1_output_port_net_x23,
      sync_out => delay0_q_net_x12
    );

  fft_stage_8_518409c227: entity work.fft_stage_8_entity_518409c227
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x14,
      in2 => reinterpret1_output_port_net_x23,
      of_in => logical1_y_net_x10,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x12,
      of_x0 => logical1_y_net_x11,
      out1 => reinterpret2_output_port_net_x15,
      out2 => reinterpret1_output_port_net_x24,
      sync_out => delay0_q_net_x13
    );

  fft_stage_9_f8166671d4: entity work.fft_stage_9_entity_f8166671d4
    port map (
      ce_1 => ce_1_sg_x501,
      clk_1 => clk_1_sg_x501,
      in1 => reinterpret2_output_port_net_x15,
      in2 => reinterpret1_output_port_net_x24,
      of_in => logical1_y_net_x11,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x13,
      of_x0 => logical1_y_net_x12,
      out1 => reinterpret2_output_port_net_x6,
      out2 => reinterpret1_output_port_net_x25,
      sync_out => delay0_q_net_x14
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core/fft_biplex_real_4x2"

entity fft_biplex_real_4x2_entity_56ec76f0c6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    pol0_in: in std_logic_vector(17 downto 0); 
    pol1_in: in std_logic_vector(17 downto 0); 
    pol2_in: in std_logic_vector(17 downto 0); 
    pol3_in: in std_logic_vector(17 downto 0); 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    pol0_out: out std_logic_vector(35 downto 0); 
    pol1_out: out std_logic_vector(35 downto 0); 
    pol2_out: out std_logic_vector(35 downto 0); 
    pol3_out: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_biplex_real_4x2_entity_56ec76f0c6;

architecture structural of fft_biplex_real_4x2_entity_56ec76f0c6 is
  signal ce_1_sg_x502: std_logic;
  signal clk_1_sg_x502: std_logic;
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal concat_y_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net_x15: std_logic;
  signal fft_shift_net_x14: std_logic_vector(31 downto 0);
  signal logical1_y_net_x14: std_logic;
  signal mux0_y_net_x3: std_logic_vector(35 downto 0);
  signal mux1_y_net_x3: std_logic_vector(35 downto 0);
  signal mux2_y_net_x3: std_logic_vector(35 downto 0);
  signal mux3_y_net_x3: std_logic_vector(35 downto 0);
  signal pol1_net_x1: std_logic_vector(17 downto 0);
  signal pol2_net_x1: std_logic_vector(17 downto 0);
  signal pol3_net_x1: std_logic_vector(17 downto 0);
  signal pol4_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x18: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x19: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x27: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x28: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x16: std_logic_vector(35 downto 0);
  signal sync_delay1_q_net_x2: std_logic;
  signal sync_net_x2: std_logic;

begin
  ce_1_sg_x502 <= ce_1;
  clk_1_sg_x502 <= clk_1;
  pol1_net_x1 <= pol0_in;
  pol2_net_x1 <= pol1_in;
  pol3_net_x1 <= pol2_in;
  pol4_net_x1 <= pol3_in;
  fft_shift_net_x14 <= shift;
  sync_net_x2 <= sync;
  of_x0 <= logical1_y_net_x14;
  pol0_out <= reinterpret1_output_port_net_x4;
  pol1_out <= reinterpret1_output_port_net_x5;
  pol2_out <= reinterpret1_output_port_net_x18;
  pol3_out <= reinterpret1_output_port_net_x19;
  sync_out <= sync_delay1_q_net_x2;

  bi_real_unscr_4x_8d809182bf: entity work.bi_real_unscr_4x_entity_8d809182bf
    port map (
      ce_1 => ce_1_sg_x502,
      clk_1 => clk_1_sg_x502,
      even => reinterpret2_output_port_net_x16,
      odd => reinterpret1_output_port_net_x27,
      sync => delay0_q_net_x15,
      pol1_out => mux0_y_net_x3,
      pol2_out => mux1_y_net_x3,
      pol3_out => mux2_y_net_x3,
      pol4_out => mux3_y_net_x3,
      sync_out => sync_delay1_q_net_x2
    );

  biplex_core_a39782552e: entity work.biplex_core_entity_a39782552e
    port map (
      ce_1 => ce_1_sg_x502,
      clk_1 => clk_1_sg_x502,
      pol1 => reinterpret1_output_port_net_x17,
      pol2 => reinterpret1_output_port_net_x28,
      shift => fft_shift_net_x14,
      sync => sync_net_x2,
      of_x0 => logical1_y_net_x14,
      out1 => reinterpret2_output_port_net_x16,
      out2 => reinterpret1_output_port_net_x27,
      sync_out => delay0_q_net_x15
    );

  even_bussify_4ef85094ca: entity work.bussify_entity_d6ea8ebb9b
    port map (
      in1 => concat_y_net_x1,
      bus_out => reinterpret1_output_port_net_x17
    );

  odd_bussify_71b77bcfac: entity work.bussify_entity_d6ea8ebb9b
    port map (
      in1 => concat_y_net_x2,
      bus_out => reinterpret1_output_port_net_x28
    );

  pol0_debus_59bc82a390: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => mux0_y_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x4
    );

  pol1_debus_f05fb45b47: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => mux1_y_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x5
    );

  pol2_debus_aaa632dab0: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => mux2_y_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x18
    );

  pol3_debus_198ff37e85: entity work.a_debus_entity_9378c272e1
    port map (
      bus_in => mux3_y_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x19
    );

  ri_to_c0_9f4b22a9bc: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => pol2_net_x1,
      re => pol1_net_x1,
      c => concat_y_net_x1
    );

  ri_to_c1_9a23b5ea50: entity work.ri_to_c_entity_7d26fbf4c5
    port map (
      im => pol4_net_x1,
      re => pol3_net_x1,
      c => concat_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_core"

entity fft_core is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_shift: in std_logic_vector(31 downto 0); 
    pol1: in std_logic_vector(17 downto 0); 
    pol2: in std_logic_vector(17 downto 0); 
    pol3: in std_logic_vector(17 downto 0); 
    pol4: in std_logic_vector(17 downto 0); 
    sync: in std_logic; 
    fft_oflow: out std_logic; 
    out_pol1: out std_logic_vector(35 downto 0); 
    out_pol2: out std_logic_vector(35 downto 0); 
    out_pol3: out std_logic_vector(35 downto 0); 
    out_pol4: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_core;

architecture structural of fft_core is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "fft_core,sysgen_core,{clock_period=10.00000000,clocking=Clock_Enables,compilation=NGC_Netlist,sample_periods=1.00000000000,testbench=0,total_blocks=9896,xilinx_adder_subtracter_block=238,xilinx_arithmetic_relational_operator_block=50,xilinx_assert_block=11,xilinx_bit_slice_extractor_block=1122,xilinx_bus_concatenator_block=385,xilinx_bus_multiplexer_block=91,xilinx_constant_block_block=464,xilinx_counter_block=65,xilinx_delay_block=309,xilinx_dual_port_random_access_memory_block=8,xilinx_gateway_in_block=6,xilinx_gateway_out_block=6,xilinx_input_scaler_block=60,xilinx_inverter_block=148,xilinx_logical_block_block=326,xilinx_multiplier_block=44,xilinx_negate_block_block=27,xilinx_register_block=22,xilinx_single_port_random_access_memory_block=24,xilinx_single_port_read_only_memory_block=6,xilinx_system_generator_block=1,xilinx_type_converter_block=96,xilinx_type_reinterpreter_block=1656,}";

  signal ce_1_sg_x503: std_logic;
  signal clk_1_sg_x503: std_logic;
  signal fft_oflow_net: std_logic;
  signal fft_shift_net: std_logic_vector(31 downto 0);
  signal out_pol1_net: std_logic_vector(35 downto 0);
  signal out_pol2_net: std_logic_vector(35 downto 0);
  signal out_pol3_net: std_logic_vector(35 downto 0);
  signal out_pol4_net: std_logic_vector(35 downto 0);
  signal pol1_net: std_logic_vector(17 downto 0);
  signal pol2_net: std_logic_vector(17 downto 0);
  signal pol3_net: std_logic_vector(17 downto 0);
  signal pol4_net: std_logic_vector(17 downto 0);
  signal sync_net: std_logic;
  signal sync_out_net: std_logic;

begin
  ce_1_sg_x503 <= ce_1;
  clk_1_sg_x503 <= clk_1;
  fft_shift_net <= fft_shift;
  pol1_net <= pol1;
  pol2_net <= pol2;
  pol3_net <= pol3;
  pol4_net <= pol4;
  sync_net <= sync;
  fft_oflow <= fft_oflow_net;
  out_pol1 <= out_pol1_net;
  out_pol2 <= out_pol2_net;
  out_pol3 <= out_pol3_net;
  out_pol4 <= out_pol4_net;
  sync_out <= sync_out_net;

  fft_biplex_real_4x2_56ec76f0c6: entity work.fft_biplex_real_4x2_entity_56ec76f0c6
    port map (
      ce_1 => ce_1_sg_x503,
      clk_1 => clk_1_sg_x503,
      pol0_in => pol1_net,
      pol1_in => pol2_net,
      pol2_in => pol3_net,
      pol3_in => pol4_net,
      shift => fft_shift_net,
      sync => sync_net,
      of_x0 => fft_oflow_net,
      pol0_out => out_pol1_net,
      pol1_out => out_pol2_net,
      pol2_out => out_pol3_net,
      pol3_out => out_pol4_net,
      sync_out => sync_out_net
    );

end structural;
