--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_a2af903969f3f923.vhd when simulating
-- the core, addsb_11_0_a2af903969f3f923. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_a2af903969f3f923 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END addsb_11_0_a2af903969f3f923;

ARCHITECTURE addsb_11_0_a2af903969f3f923_a OF addsb_11_0_a2af903969f3f923 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_a2af903969f3f923
  PORT (
    a : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_a2af903969f3f923 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 12,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000",
      c_b_width => 12,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 12,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_a2af903969f3f923
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_a2af903969f3f923_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_efdf1b1b05926829.vhd when simulating
-- the core, dmg_72_efdf1b1b05926829. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_efdf1b1b05926829 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_efdf1b1b05926829;

ARCHITECTURE dmg_72_efdf1b1b05926829_a OF dmg_72_efdf1b1b05926829 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_efdf1b1b05926829
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_efdf1b1b05926829 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_efdf1b1b05926829.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_efdf1b1b05926829
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_efdf1b1b05926829_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_9f585cf1e3329833.vhd when simulating
-- the core, bmg_72_9f585cf1e3329833. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_9f585cf1e3329833 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_9f585cf1e3329833;

ARCHITECTURE bmg_72_9f585cf1e3329833_a OF bmg_72_9f585cf1e3329833 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_9f585cf1e3329833
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_9f585cf1e3329833 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 10,
      c_addrb_width => 10,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_9f585cf1e3329833.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 1024,
      c_read_depth_b => 1024,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 1024,
      c_write_depth_b => 1024,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_9f585cf1e3329833
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_9f585cf1e3329833_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_618ffcc3f0781f68.vhd when simulating
-- the core, bmg_72_618ffcc3f0781f68. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_618ffcc3f0781f68 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_618ffcc3f0781f68;

ARCHITECTURE bmg_72_618ffcc3f0781f68_a OF bmg_72_618ffcc3f0781f68 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_618ffcc3f0781f68
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_618ffcc3f0781f68 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 8,
      c_addrb_width => 8,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_618ffcc3f0781f68.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 5,
      c_read_depth_a => 256,
      c_read_depth_b => 256,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 256,
      c_write_depth_b => 256,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_618ffcc3f0781f68
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_618ffcc3f0781f68_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_15a84ff1ccdd3419.vhd when simulating
-- the core, bmg_72_15a84ff1ccdd3419. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_15a84ff1ccdd3419 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_15a84ff1ccdd3419;

ARCHITECTURE bmg_72_15a84ff1ccdd3419_a OF bmg_72_15a84ff1ccdd3419 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_15a84ff1ccdd3419
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_15a84ff1ccdd3419 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 10,
      c_addrb_width => 10,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_15a84ff1ccdd3419.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 1024,
      c_read_depth_b => 1024,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 1024,
      c_write_depth_b => 1024,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_15a84ff1ccdd3419
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_15a84ff1ccdd3419_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_47829d325bbb998a.vhd when simulating
-- the core, addsb_11_0_47829d325bbb998a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_47829d325bbb998a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END addsb_11_0_47829d325bbb998a;

ARCHITECTURE addsb_11_0_47829d325bbb998a_a OF addsb_11_0_47829d325bbb998a IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_47829d325bbb998a
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_47829d325bbb998a USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 13,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000",
      c_b_width => 13,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 13,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_47829d325bbb998a
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_47829d325bbb998a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_a0497faccc62b6b2.vhd when simulating
-- the core, addsb_11_0_a0497faccc62b6b2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_a0497faccc62b6b2 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END addsb_11_0_a0497faccc62b6b2;

ARCHITECTURE addsb_11_0_a0497faccc62b6b2_a OF addsb_11_0_a0497faccc62b6b2 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_a0497faccc62b6b2
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_a0497faccc62b6b2 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 20,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000",
      c_b_width => 20,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 20,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_a0497faccc62b6b2
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_a0497faccc62b6b2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_5ed93725c6f3d1db.vhd when simulating
-- the core, bmg_72_5ed93725c6f3d1db. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_5ed93725c6f3d1db IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_5ed93725c6f3d1db;

ARCHITECTURE bmg_72_5ed93725c6f3d1db_a OF bmg_72_5ed93725c6f3d1db IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_5ed93725c6f3d1db
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_5ed93725c6f3d1db USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_5ed93725c6f3d1db.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 5,
      c_read_depth_a => 64,
      c_read_depth_b => 64,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 64,
      c_write_depth_b => 64,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_5ed93725c6f3d1db
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_5ed93725c6f3d1db_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_59920783799a8e86.vhd when simulating
-- the core, addsb_11_0_59920783799a8e86. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_59920783799a8e86 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_59920783799a8e86;

ARCHITECTURE addsb_11_0_59920783799a8e86_a OF addsb_11_0_59920783799a8e86 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_59920783799a8e86
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_59920783799a8e86 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_59920783799a8e86
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_59920783799a8e86_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_180432cd81ea5a8d.vhd when simulating
-- the core, bmg_72_180432cd81ea5a8d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_180432cd81ea5a8d IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END bmg_72_180432cd81ea5a8d;

ARCHITECTURE bmg_72_180432cd81ea5a8d_a OF bmg_72_180432cd81ea5a8d IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_180432cd81ea5a8d
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_180432cd81ea5a8d USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_180432cd81ea5a8d.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 2,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 12,
      c_read_width_b => 12,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 12,
      c_write_width_b => 12,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_180432cd81ea5a8d
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_180432cd81ea5a8d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_7eed1f270da26adb.vhd when simulating
-- the core, bmg_72_7eed1f270da26adb. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_7eed1f270da26adb IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END bmg_72_7eed1f270da26adb;

ARCHITECTURE bmg_72_7eed1f270da26adb_a OF bmg_72_7eed1f270da26adb IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_7eed1f270da26adb
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_7eed1f270da26adb USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 11,
      c_addrb_width => 11,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_7eed1f270da26adb.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 3,
      c_read_depth_a => 2048,
      c_read_depth_b => 2048,
      c_read_width_a => 9,
      c_read_width_b => 9,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 2048,
      c_write_depth_b => 2048,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 9,
      c_write_width_b => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_7eed1f270da26adb
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_7eed1f270da26adb_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_fa6496d84f038019.vhd when simulating
-- the core, bmg_72_fa6496d84f038019. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_fa6496d84f038019 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END bmg_72_fa6496d84f038019;

ARCHITECTURE bmg_72_fa6496d84f038019_a OF bmg_72_fa6496d84f038019 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_fa6496d84f038019
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_fa6496d84f038019 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_fa6496d84f038019.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 2,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 4,
      c_read_width_b => 4,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 4,
      c_write_width_b => 4,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_fa6496d84f038019
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_fa6496d84f038019_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_80a4fb0fcb4866f6.vhd when simulating
-- the core, addsb_11_0_80a4fb0fcb4866f6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_80a4fb0fcb4866f6 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END addsb_11_0_80a4fb0fcb4866f6;

ARCHITECTURE addsb_11_0_80a4fb0fcb4866f6_a OF addsb_11_0_80a4fb0fcb4866f6 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_80a4fb0fcb4866f6
  PORT (
    a : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_80a4fb0fcb4866f6 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 22,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000000",
      c_b_width => 22,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 22,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_80a4fb0fcb4866f6
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_80a4fb0fcb4866f6_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_3d733db2a81768b0.vhd when simulating
-- the core, bmg_72_3d733db2a81768b0. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_3d733db2a81768b0 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_3d733db2a81768b0;

ARCHITECTURE bmg_72_3d733db2a81768b0_a OF bmg_72_3d733db2a81768b0 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_3d733db2a81768b0
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_3d733db2a81768b0 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 7,
      c_addrb_width => 7,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_3d733db2a81768b0.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 5,
      c_read_depth_a => 128,
      c_read_depth_b => 128,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 128,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_3d733db2a81768b0
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_3d733db2a81768b0_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_1c323e86177437db.vhd when simulating
-- the core, dmg_72_1c323e86177437db. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_1c323e86177437db IS
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_1c323e86177437db;

ARCHITECTURE dmg_72_1c323e86177437db_a OF dmg_72_1c323e86177437db IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_1c323e86177437db
  PORT (
    a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_1c323e86177437db USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 5,
      c_default_data => "0",
      c_depth => 32,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_1c323e86177437db.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_1c323e86177437db
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_1c323e86177437db_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_18f6f1cec46d694e.vhd when simulating
-- the core, addsb_11_0_18f6f1cec46d694e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_18f6f1cec46d694e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_18f6f1cec46d694e;

ARCHITECTURE addsb_11_0_18f6f1cec46d694e_a OF addsb_11_0_18f6f1cec46d694e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_18f6f1cec46d694e
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_18f6f1cec46d694e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_18f6f1cec46d694e
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_18f6f1cec46d694e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_ce7e9961dfcc2802.vhd when simulating
-- the core, bmg_72_ce7e9961dfcc2802. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_ce7e9961dfcc2802 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END bmg_72_ce7e9961dfcc2802;

ARCHITECTURE bmg_72_ce7e9961dfcc2802_a OF bmg_72_ce7e9961dfcc2802 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_ce7e9961dfcc2802
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_ce7e9961dfcc2802 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_ce7e9961dfcc2802.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 2,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 12,
      c_read_width_b => 12,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 12,
      c_write_width_b => 12,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_ce7e9961dfcc2802
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_ce7e9961dfcc2802_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_8574240a262aac9a.vhd when simulating
-- the core, bmg_72_8574240a262aac9a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_8574240a262aac9a IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END bmg_72_8574240a262aac9a;

ARCHITECTURE bmg_72_8574240a262aac9a_a OF bmg_72_8574240a262aac9a IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_8574240a262aac9a
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_8574240a262aac9a USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_8574240a262aac9a.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 2,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 12,
      c_read_width_b => 12,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 12,
      c_write_width_b => 12,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_8574240a262aac9a
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_8574240a262aac9a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_e02664f04ec6e0c0.vhd when simulating
-- the core, bmg_72_e02664f04ec6e0c0. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_e02664f04ec6e0c0 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_e02664f04ec6e0c0;

ARCHITECTURE bmg_72_e02664f04ec6e0c0_a OF bmg_72_e02664f04ec6e0c0 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_e02664f04ec6e0c0
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_e02664f04ec6e0c0 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 9,
      c_addrb_width => 9,
      c_algorithm => 0,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_e02664f04ec6e0c0.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 5,
      c_read_depth_a => 512,
      c_read_depth_b => 512,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 512,
      c_write_depth_b => 512,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_e02664f04ec6e0c0
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_e02664f04ec6e0c0_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_c055560701350b3e.vhd when simulating
-- the core, addsb_11_0_c055560701350b3e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_c055560701350b3e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END addsb_11_0_c055560701350b3e;

ARCHITECTURE addsb_11_0_c055560701350b3e_a OF addsb_11_0_c055560701350b3e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_c055560701350b3e
  PORT (
    a : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_c055560701350b3e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 22,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000000",
      c_b_width => 22,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 22,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_c055560701350b3e
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_c055560701350b3e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_6e641a09b813308f.vhd when simulating
-- the core, addsb_11_0_6e641a09b813308f. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_6e641a09b813308f IS
  PORT (
    a : IN STD_LOGIC_VECTOR(38 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(38 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(38 DOWNTO 0)
  );
END addsb_11_0_6e641a09b813308f;

ARCHITECTURE addsb_11_0_6e641a09b813308f_a OF addsb_11_0_6e641a09b813308f IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_6e641a09b813308f
  PORT (
    a : IN STD_LOGIC_VECTOR(38 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(38 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(38 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_6e641a09b813308f USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 39,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000000000000000000000000",
      c_b_width => 39,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 39,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_6e641a09b813308f
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_6e641a09b813308f_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_9d950569c0d7f9e8.vhd when simulating
-- the core, bmg_72_9d950569c0d7f9e8. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_9d950569c0d7f9e8 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END bmg_72_9d950569c0d7f9e8;

ARCHITECTURE bmg_72_9d950569c0d7f9e8_a OF bmg_72_9d950569c0d7f9e8 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_9d950569c0d7f9e8
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_9d950569c0d7f9e8 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 11,
      c_addrb_width => 11,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 1,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_9d950569c0d7f9e8.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 2048,
      c_read_depth_b => 2048,
      c_read_width_a => 18,
      c_read_width_b => 18,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 2048,
      c_write_depth_b => 2048,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 18,
      c_write_width_b => 18,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_9d950569c0d7f9e8
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_9d950569c0d7f9e8_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_ff0037ba5117ccc6.vhd when simulating
-- the core, addsb_11_0_ff0037ba5117ccc6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_ff0037ba5117ccc6 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
  );
END addsb_11_0_ff0037ba5117ccc6;

ARCHITECTURE addsb_11_0_ff0037ba5117ccc6_a OF addsb_11_0_ff0037ba5117ccc6 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_ff0037ba5117ccc6
  PORT (
    a : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_ff0037ba5117ccc6 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 21,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000000",
      c_b_width => 21,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 21,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_ff0037ba5117ccc6
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_ff0037ba5117ccc6_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_0b9daa5d24360c6e.vhd when simulating
-- the core, addsb_11_0_0b9daa5d24360c6e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_0b9daa5d24360c6e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_0b9daa5d24360c6e;

ARCHITECTURE addsb_11_0_0b9daa5d24360c6e_a OF addsb_11_0_0b9daa5d24360c6e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_0b9daa5d24360c6e
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_0b9daa5d24360c6e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_0b9daa5d24360c6e
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_0b9daa5d24360c6e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_d20b02a9f8239c7a.vhd when simulating
-- the core, dmg_72_d20b02a9f8239c7a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_d20b02a9f8239c7a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_d20b02a9f8239c7a;

ARCHITECTURE dmg_72_d20b02a9f8239c7a_a OF dmg_72_d20b02a9f8239c7a IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_d20b02a9f8239c7a
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_d20b02a9f8239c7a USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_d20b02a9f8239c7a.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_d20b02a9f8239c7a
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_d20b02a9f8239c7a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_505931c5b3ea228e.vhd when simulating
-- the core, dmg_72_505931c5b3ea228e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_505931c5b3ea228e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END dmg_72_505931c5b3ea228e;

ARCHITECTURE dmg_72_505931c5b3ea228e_a OF dmg_72_505931c5b3ea228e IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_505931c5b3ea228e
  PORT (
    a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    d : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpra : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    clk : IN STD_LOGIC;
    we : IN STD_LOGIC;
    spo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
    dpo : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_505931c5b3ea228e USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 4,
      c_default_data => "0",
      c_depth => 16,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 1,
      c_has_dpo => 1,
      c_has_dpra => 1,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 1,
      c_mem_init_file => "dmg_72_505931c5b3ea228e.mif",
      c_mem_type => 2,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 18
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_505931c5b3ea228e
  PORT MAP (
    a => a,
    d => d,
    dpra => dpra,
    clk => clk,
    we => we,
    spo => spo,
    dpo => dpo
  );
-- synthesis translate_on

END dmg_72_505931c5b3ea228e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_3af1276811d12ede.vhd when simulating
-- the core, addsb_11_0_3af1276811d12ede. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_3af1276811d12ede IS
  PORT (
    a : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
  );
END addsb_11_0_3af1276811d12ede;

ARCHITECTURE addsb_11_0_3af1276811d12ede_a OF addsb_11_0_3af1276811d12ede IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_3af1276811d12ede
  PORT (
    a : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(20 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(20 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_3af1276811d12ede USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 21,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000000",
      c_b_width => 21,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 21,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_3af1276811d12ede
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_3af1276811d12ede_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_6bbb8fb0d8f20abe.vhd when simulating
-- the core, addsb_11_0_6bbb8fb0d8f20abe. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_6bbb8fb0d8f20abe IS
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END addsb_11_0_6bbb8fb0d8f20abe;

ARCHITECTURE addsb_11_0_6bbb8fb0d8f20abe_a OF addsb_11_0_6bbb8fb0d8f20abe IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_6bbb8fb0d8f20abe
  PORT (
    a : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_6bbb8fb0d8f20abe USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 20,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000",
      c_b_width => 20,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 20,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_6bbb8fb0d8f20abe
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_6bbb8fb0d8f20abe_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_c9b173d075a3b6d7.vhd when simulating
-- the core, addsb_11_0_c9b173d075a3b6d7. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_c9b173d075a3b6d7 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END addsb_11_0_c9b173d075a3b6d7;

ARCHITECTURE addsb_11_0_c9b173d075a3b6d7_a OF addsb_11_0_c9b173d075a3b6d7 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_c9b173d075a3b6d7
  PORT (
    a : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(18 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(18 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_c9b173d075a3b6d7 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 19,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000",
      c_b_width => 19,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 1,
      c_latency => 1,
      c_out_width => 19,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_c9b173d075a3b6d7
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_c9b173d075a3b6d7_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_77dc1780892a0930.vhd when simulating
-- the core, bmg_72_77dc1780892a0930. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_77dc1780892a0930 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END bmg_72_77dc1780892a0930;

ARCHITECTURE bmg_72_77dc1780892a0930_a OF bmg_72_77dc1780892a0930 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_77dc1780892a0930
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(35 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(35 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_77dc1780892a0930 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 12,
      c_addrb_width => 12,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 1,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_77dc1780892a0930.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 0,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 4096,
      c_read_depth_b => 4096,
      c_read_width_a => 36,
      c_read_width_b => 36,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 4096,
      c_write_depth_b => 4096,
      c_write_mode_a => "READ_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 36,
      c_write_width_b => 36,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_77dc1780892a0930
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_77dc1780892a0930_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2016 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_1f22b9fac024cf00.vhd when simulating
-- the core, addsb_11_0_1f22b9fac024cf00. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_1f22b9fac024cf00 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(22 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(22 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(22 DOWNTO 0)
  );
END addsb_11_0_1f22b9fac024cf00;

ARCHITECTURE addsb_11_0_1f22b9fac024cf00_a OF addsb_11_0_1f22b9fac024cf00 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_1f22b9fac024cf00
  PORT (
    a : IN STD_LOGIC_VECTOR(22 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(22 DOWNTO 0);
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    s : OUT STD_LOGIC_VECTOR(22 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_1f22b9fac024cf00 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 23,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000000",
      c_b_width => 23,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 1,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 1,
      c_out_width => 23,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_1f22b9fac024cf00
  PORT MAP (
    a => a,
    b => b,
    clk => clk,
    ce => ce,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_1f22b9fac024cf00_a;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_e110f0a1fc is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_e110f0a1fc;


architecture behavior of counter_e110f0a1fc is
  signal count_reg_20_23: unsigned((12 - 1) downto 0) := "000000000000";
  signal count_reg_20_23_rst: std_logic;
  signal rel_34_8: boolean;
  signal rst_limit_join_34_5: boolean;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((13 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  rel_34_8 <= count_reg_20_23 = std_logic_vector_to_unsigned("111111111100");
  proc_if_34_5: process (rel_34_8)
  is
  begin
    if rel_34_8 then
      rst_limit_join_34_5 <= true;
    else 
      rst_limit_join_34_5 <= false;
    end if;
  end process proc_if_34_5;
  bool_44_4 <= false or rst_limit_join_34_5;
  proc_if_44_1: process (bool_44_4, count_reg_20_23, rst_limit_join_34_5)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= rst_limit_join_34_5;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlspram_fft_astro_devel_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
    );
  port (
    data_in: in std_logic_vector(c_width - 1 downto 0);
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    we: in std_logic_vector(0 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data_out: out std_logic_vector(c_width - 1 downto 0)
  );
end xlspram_fft_astro_devel_core ;
architecture behavior of xlspram_fft_astro_devel_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_data_out, dly_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_we, core_ce, sinit: std_logic;
  component bmg_72_77dc1780892a0930
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_77dc1780892a0930:
    component is true;
  attribute fpga_dont_touch of bmg_72_77dc1780892a0930:
    component is "true";
  attribute box_type of bmg_72_77dc1780892a0930:
    component  is "black_box";
  component bmg_72_fa6496d84f038019
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_fa6496d84f038019:
    component is true;
  attribute fpga_dont_touch of bmg_72_fa6496d84f038019:
    component is "true";
  attribute box_type of bmg_72_fa6496d84f038019:
    component  is "black_box";
  component bmg_72_7eed1f270da26adb
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      dina: in std_logic_vector(c_width - 1 downto 0);
      wea: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_7eed1f270da26adb:
    component is true;
  attribute fpga_dont_touch of bmg_72_7eed1f270da26adb:
    component is "true";
  attribute box_type of bmg_72_7eed1f270da26adb:
    component  is "black_box";
begin
  data_out <= dly_data_out;
  core_we <= we(0);
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_77dc1780892a0930")) generate
    core_instance0: bmg_72_77dc1780892a0930
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_fa6496d84f038019")) generate
    core_instance1: bmg_72_fa6496d84f038019
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  comp2: if ((core_name0 = "bmg_72_7eed1f270da26adb")) generate
    core_instance2: bmg_72_7eed1f270da26adb
      port map (
                                        addra => addr,
        clka => clk,
        dina => data_in,
        wea(0) => core_we,
        ena => core_ce,
        douta => core_data_out
      );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => dly_data_out
      );
  end generate;
  latency_1: if (latency <= 1) generate
    dly_data_out <= core_data_out;
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9a0fa0f632 is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9a0fa0f632;


architecture behavior of reinterpret_9a0fa0f632 is
  signal input_port_1_40: unsigned((18 - 1) downto 0);
  signal output_port_5_5_force: signed((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlslice is
    generic (
        new_msb      : integer := 9;
        new_lsb      : integer := 1;
        x_width      : integer := 16;
        y_width      : integer := 8);
    port (
        x : in std_logic_vector (x_width-1 downto 0);
        y : out std_logic_vector (y_width-1 downto 0));
end xlslice;
architecture behavior of xlslice is
begin
    y <= x(new_msb downto new_lsb);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_bc4405cd1e is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_bc4405cd1e;


architecture behavior of reinterpret_bc4405cd1e is
  signal input_port_1_40: signed((19 - 1) downto 0);
  signal output_port_5_5_force: unsigned((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub_fft_astro_devel_core is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub_fft_astro_devel_core;
architecture behavior of xladdsub_fft_astro_devel_core is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_59920783799a8e86
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_ff0037ba5117ccc6
    port (
          a: in std_logic_vector(21 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(21 - 1 downto 0)
    );
  end component;
  component addsb_11_0_18f6f1cec46d694e
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_0b9daa5d24360c6e
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_80a4fb0fcb4866f6
    port (
          a: in std_logic_vector(22 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(22 - 1 downto 0)
    );
  end component;
  component addsb_11_0_3af1276811d12ede
    port (
          a: in std_logic_vector(21 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(21 - 1 downto 0)
    );
  end component;
  component addsb_11_0_c9b173d075a3b6d7
    port (
          a: in std_logic_vector(19 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(19 - 1 downto 0)
    );
  end component;
  component addsb_11_0_6bbb8fb0d8f20abe
    port (
          a: in std_logic_vector(20 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(20 - 1 downto 0)
    );
  end component;
  component addsb_11_0_1f22b9fac024cf00
    port (
          a: in std_logic_vector(23 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(23 - 1 downto 0)
    );
  end component;
  component addsb_11_0_c055560701350b3e
    port (
          a: in std_logic_vector(22 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(22 - 1 downto 0)
    );
  end component;
  component addsb_11_0_a0497faccc62b6b2
    port (
          a: in std_logic_vector(20 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(20 - 1 downto 0)
    );
  end component;
  component addsb_11_0_6e641a09b813308f
    port (
          a: in std_logic_vector(39 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(39 - 1 downto 0)
    );
  end component;
  component addsb_11_0_a2af903969f3f923
    port (
          a: in std_logic_vector(12 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(12 - 1 downto 0)
    );
  end component;
  component addsb_11_0_47829d325bbb998a
    port (
          a: in std_logic_vector(13 - 1 downto 0);
    clk: in std_logic:= '0';
    ce: in std_logic:= '0';
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(13 - 1 downto 0)
    );
  end component;
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_59920783799a8e86")) generate
    core_instance0: addsb_11_0_59920783799a8e86
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp1: if ((core_name0 = "addsb_11_0_ff0037ba5117ccc6")) generate
    core_instance1: addsb_11_0_ff0037ba5117ccc6
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_18f6f1cec46d694e")) generate
    core_instance2: addsb_11_0_18f6f1cec46d694e
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp3: if ((core_name0 = "addsb_11_0_0b9daa5d24360c6e")) generate
    core_instance3: addsb_11_0_0b9daa5d24360c6e
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp4: if ((core_name0 = "addsb_11_0_80a4fb0fcb4866f6")) generate
    core_instance4: addsb_11_0_80a4fb0fcb4866f6
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp5: if ((core_name0 = "addsb_11_0_3af1276811d12ede")) generate
    core_instance5: addsb_11_0_3af1276811d12ede
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp6: if ((core_name0 = "addsb_11_0_c9b173d075a3b6d7")) generate
    core_instance6: addsb_11_0_c9b173d075a3b6d7
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp7: if ((core_name0 = "addsb_11_0_6bbb8fb0d8f20abe")) generate
    core_instance7: addsb_11_0_6bbb8fb0d8f20abe
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp8: if ((core_name0 = "addsb_11_0_1f22b9fac024cf00")) generate
    core_instance8: addsb_11_0_1f22b9fac024cf00
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp9: if ((core_name0 = "addsb_11_0_c055560701350b3e")) generate
    core_instance9: addsb_11_0_c055560701350b3e
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp10: if ((core_name0 = "addsb_11_0_a0497faccc62b6b2")) generate
    core_instance10: addsb_11_0_a0497faccc62b6b2
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp11: if ((core_name0 = "addsb_11_0_6e641a09b813308f")) generate
    core_instance11: addsb_11_0_6e641a09b813308f
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp12: if ((core_name0 = "addsb_11_0_a2af903969f3f923")) generate
    core_instance12: addsb_11_0_a2af903969f3f923
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  comp13: if ((core_name0 = "addsb_11_0_47829d325bbb998a")) generate
    core_instance13: addsb_11_0_47829d325bbb998a
      port map (
         a => full_a,
         clk => clk,
         ce => internal_ce,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a246e373e7 is
  port (
    in0 : in std_logic_vector((18 - 1) downto 0);
    in1 : in std_logic_vector((18 - 1) downto 0);
    in2 : in std_logic_vector((18 - 1) downto 0);
    in3 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((72 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a246e373e7;


architecture behavior of concat_a246e373e7 is
  signal in0_1_23: unsigned((18 - 1) downto 0);
  signal in1_1_27: unsigned((18 - 1) downto 0);
  signal in2_1_31: unsigned((18 - 1) downto 0);
  signal in3_1_35: unsigned((18 - 1) downto 0);
  signal y_2_1_concat: unsigned((72 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_580feec131 is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_580feec131;


architecture behavior of reinterpret_580feec131 is
  signal input_port_1_40: signed((18 - 1) downto 0);
  signal output_port_5_5_force: unsigned((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_504cae28bd is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_504cae28bd;


architecture behavior of concat_504cae28bd is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((20 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4709ea49b5 is
  port (
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4709ea49b5;


architecture behavior of constant_4709ea49b5 is
begin
  op <= "0000000000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_f661f8d9b7 is
  port (
    input_port : in std_logic_vector((20 - 1) downto 0);
    output_port : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_f661f8d9b7;


architecture behavior of reinterpret_f661f8d9b7 is
  signal input_port_1_40: unsigned((20 - 1) downto 0);
  signal output_port_5_5_force: signed((20 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d2180c9169 is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d2180c9169;


architecture behavior of reinterpret_d2180c9169 is
  signal input_port_1_40: unsigned((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_938d99ac11 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_938d99ac11;


architecture behavior of logical_938d99ac11 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_63700884f5 is
  port (
    input_port : in std_logic_vector((19 - 1) downto 0);
    output_port : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_63700884f5;


architecture behavior of reinterpret_63700884f5 is
  signal input_port_1_40: unsigned((19 - 1) downto 0);
  signal output_port_5_5_force: signed((19 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9306b5127f is
  port (
    input_port : in std_logic_vector((18 - 1) downto 0);
    output_port : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9306b5127f;


architecture behavior of reinterpret_9306b5127f is
  signal input_port_1_40: unsigned((18 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2aea51ccde is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((19 - 1) downto 0);
    in2 : in std_logic_vector((19 - 1) downto 0);
    in3 : in std_logic_vector((19 - 1) downto 0);
    y : out std_logic_vector((76 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2aea51ccde;


architecture behavior of concat_2aea51ccde is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((19 - 1) downto 0);
  signal in2_1_31: unsigned((19 - 1) downto 0);
  signal in3_1_35: unsigned((19 - 1) downto 0);
  signal y_2_1_concat: unsigned((76 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity scale_9f61027ba4 is
  port (
    ip : in std_logic_vector((19 - 1) downto 0);
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end scale_9f61027ba4;


architecture behavior of scale_9f61027ba4 is
  signal ip_17_23: signed((19 - 1) downto 0);
begin
  ip_17_23 <= std_logic_vector_to_signed(ip);
  op <= signed_to_std_logic_vector(ip_17_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_b198bd62b0 is
  port (
    in0 : in std_logic_vector((18 - 1) downto 0);
    in1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_b198bd62b0;


architecture behavior of concat_b198bd62b0 is
  signal in0_1_23: unsigned((18 - 1) downto 0);
  signal in1_1_27: unsigned((18 - 1) downto 0);
  signal y_2_1_concat: unsigned((36 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_86b044698f is
  port (
    input_port : in std_logic_vector((36 - 1) downto 0);
    output_port : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_86b044698f;


architecture behavior of reinterpret_86b044698f is
  signal input_port_1_40: unsigned((36 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_f983e30a8b is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_f983e30a8b;


architecture behavior of negate_f983e30a8b is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (1 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    0 => "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal cast_internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(0);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  cast_internal_ip_40_3_convert <= s2s_cast(internal_ip_join_30_1, 17, 18, 17);
  op_mem_48_20_push_front_pop_back_en <= '0';
  op <= signed_to_std_logic_vector(cast_internal_ip_40_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_6699ee0916 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_6699ee0916;


architecture behavior of delay_6699ee0916 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_81130c7f2d is
  port (
    input_port : in std_logic_vector((1 - 1) downto 0);
    output_port : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_81130c7f2d;


architecture behavior of reinterpret_81130c7f2d is
  signal input_port_1_40: unsigned((1 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4bb6f691f7 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((36 - 1) downto 0);
    d1 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4bb6f691f7;


architecture behavior of mux_4bb6f691f7 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((36 - 1) downto 0);
  signal d1_1_27: std_logic_vector((36 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((36 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_112d91c147 is
  port (
    input_port : in std_logic_vector((1 - 1) downto 0);
    output_port : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_112d91c147;


architecture behavior of reinterpret_112d91c147 is
  signal input_port_1_40: boolean;
  signal output_port_7_5_convert: unsigned((1 - 1) downto 0);
begin
  input_port_1_40 <= ((input_port) = "1");
  output_port_7_5_convert <= u2u_cast(std_logic_vector_to_unsigned(boolean_to_vector(input_port_1_40)), 0, 1, 0);
  output_port <= unsigned_to_std_logic_vector(output_port_7_5_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e055964d40 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e055964d40;


architecture behavior of delay_e055964d40 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (13 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(12);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 12 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_c48d6dcab5 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_c48d6dcab5;


architecture behavior of counter_c48d6dcab5 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((13 - 1) downto 0) := "0000000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((14 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0000000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("0000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e47f8076b8 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e47f8076b8;


architecture behavior of constant_e47f8076b8 is
begin
  op <= "1000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_54e7975215 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54e7975215;


architecture behavior of relational_54e7975215 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_9f02caa990 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_9f02caa990;


architecture behavior of delay_9f02caa990 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_6096a10519 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_6096a10519;


architecture behavior of delay_6096a10519 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (13 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(12);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 12 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_75275f6c4a is
  port (
    input_port : in std_logic_vector((12 - 1) downto 0);
    output_port : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_75275f6c4a;


architecture behavior of reinterpret_75275f6c4a is
  signal input_port_1_40: unsigned((12 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d610556e85 is
  port (
    input_port : in std_logic_vector((4 - 1) downto 0);
    output_port : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d610556e85;


architecture behavior of reinterpret_d610556e85 is
  signal input_port_1_40: unsigned((4 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e4837c85a3 is
  port (
    in0 : in std_logic_vector((4 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    in2 : in std_logic_vector((4 - 1) downto 0);
    in3 : in std_logic_vector((4 - 1) downto 0);
    in4 : in std_logic_vector((4 - 1) downto 0);
    in5 : in std_logic_vector((4 - 1) downto 0);
    in6 : in std_logic_vector((4 - 1) downto 0);
    in7 : in std_logic_vector((4 - 1) downto 0);
    in8 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e4837c85a3;


architecture behavior of concat_e4837c85a3 is
  signal in0_1_23: unsigned((4 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal in2_1_31: unsigned((4 - 1) downto 0);
  signal in3_1_35: unsigned((4 - 1) downto 0);
  signal in4_1_39: unsigned((4 - 1) downto 0);
  signal in5_1_43: unsigned((4 - 1) downto 0);
  signal in6_1_47: unsigned((4 - 1) downto 0);
  signal in7_1_51: unsigned((4 - 1) downto 0);
  signal in8_1_55: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((36 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_336ab7141a is
  port (
    in0 : in std_logic_vector((12 - 1) downto 0);
    in1 : in std_logic_vector((12 - 1) downto 0);
    in2 : in std_logic_vector((12 - 1) downto 0);
    in3 : in std_logic_vector((12 - 1) downto 0);
    in4 : in std_logic_vector((12 - 1) downto 0);
    in5 : in std_logic_vector((12 - 1) downto 0);
    in6 : in std_logic_vector((12 - 1) downto 0);
    in7 : in std_logic_vector((12 - 1) downto 0);
    in8 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((108 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_336ab7141a;


architecture behavior of concat_336ab7141a is
  signal in0_1_23: unsigned((12 - 1) downto 0);
  signal in1_1_27: unsigned((12 - 1) downto 0);
  signal in2_1_31: unsigned((12 - 1) downto 0);
  signal in3_1_35: unsigned((12 - 1) downto 0);
  signal in4_1_39: unsigned((12 - 1) downto 0);
  signal in5_1_43: unsigned((12 - 1) downto 0);
  signal in6_1_47: unsigned((12 - 1) downto 0);
  signal in7_1_51: unsigned((12 - 1) downto 0);
  signal in8_1_55: unsigned((12 - 1) downto 0);
  signal y_2_1_concat: unsigned((108 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer :=  0;
           reset        : integer :=  0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        rst     : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if ((reg_retiming = 0) and (reset = 0)) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if ((reg_retiming = 1) or (reset = 1)) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => rst,
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_0cc72cd991 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_0cc72cd991;


architecture behavior of concat_0cc72cd991 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_bdaf6c9e55 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_bdaf6c9e55;


architecture behavior of delay_bdaf6c9e55 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (4 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(3);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_50be3b5040 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_50be3b5040;


architecture behavior of constant_50be3b5040 is
begin
  op <= "0000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0c8736a503 is
  port (
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0c8736a503;


architecture behavior of constant_0c8736a503 is
begin
  op <= "0000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_eb4d9e2dad is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((13 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_eb4d9e2dad;


architecture behavior of counter_eb4d9e2dad is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((13 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((13 - 1) downto 0);
  signal count_reg_20_23: unsigned((13 - 1) downto 0) := "0000000000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((15 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((15 - 1) downto 0);
  signal count_reg_join_48_3: signed((15 - 1) downto 0);
  signal count_reg_join_44_1: signed((15 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((13 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 15, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("000000000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 15, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 13, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_80f90b97d0 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_80f90b97d0;


architecture behavior of logical_80f90b97d0 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1bef4ba0e4 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1bef4ba0e4;


architecture behavior of mux_1bef4ba0e4 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal unregy_join_6_1: std_logic;
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= std_logic_to_vector(unregy_join_6_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6dfa374756 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6dfa374756;


architecture behavior of relational_6dfa374756 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2550da35d2 is
  port (
    a : in std_logic_vector((13 - 1) downto 0);
    b : in std_logic_vector((13 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2550da35d2;


architecture behavior of relational_2550da35d2 is
  signal a_1_31: unsigned((13 - 1) downto 0);
  signal b_1_34: unsigned((13 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_c53de546ea is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_c53de546ea;


architecture behavior of delay_c53de546ea is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (4 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(3);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_fa260f7d22 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_fa260f7d22;


architecture behavior of delay_fa260f7d22 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (7 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(6);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 6 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_486acbf0b9 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_486acbf0b9;


architecture behavior of counter_486acbf0b9 is
  signal rst_1_40: boolean;
  signal en_1_45: boolean;
  signal count_reg_20_23: unsigned((13 - 1) downto 0) := "0000000000000";
  signal count_reg_20_23_rst: std_logic;
  signal count_reg_20_23_en: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((14 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0000000000000";
      elsif ((ce = '1') and (count_reg_20_23_en = '1')) then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("0000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23, en_1_45)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    elsif en_1_45 then
      count_reg_join_44_1_rst <= '0';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    elsif en_1_45 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_85c2ef968b is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_85c2ef968b;


architecture behavior of delay_85c2ef968b is
  signal d_1_22: std_logic_vector((1 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0",
    "0",
    "0");
  signal op_mem_20_24_front_din: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_b1290993d1 is
  port (
    d : in std_logic_vector((12 - 1) downto 0);
    q : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_b1290993d1;


architecture behavior of delay_b1290993d1 is
  signal d_1_22: std_logic_vector((12 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000",
    "000000000000",
    "000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_25f2d74a2a is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_25f2d74a2a;


architecture behavior of mux_25f2d74a2a is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000");
  signal pipe_16_22_front_din: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_fft_astro_devel_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_fft_astro_devel_core ;
architecture behavior of xlsprom_fft_astro_devel_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_ce, sinit: std_logic;
  component bmg_72_180432cd81ea5a8d
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_180432cd81ea5a8d:
    component is true;
  attribute fpga_dont_touch of bmg_72_180432cd81ea5a8d:
    component is "true";
  attribute box_type of bmg_72_180432cd81ea5a8d:
    component  is "black_box";
  component bmg_72_8574240a262aac9a
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_8574240a262aac9a:
    component is true;
  attribute fpga_dont_touch of bmg_72_8574240a262aac9a:
    component is "true";
  attribute box_type of bmg_72_8574240a262aac9a:
    component  is "black_box";
  component bmg_72_ce7e9961dfcc2802
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_ce7e9961dfcc2802:
    component is true;
  attribute fpga_dont_touch of bmg_72_ce7e9961dfcc2802:
    component is "true";
  attribute box_type of bmg_72_ce7e9961dfcc2802:
    component  is "black_box";
  component bmg_72_e02664f04ec6e0c0
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_e02664f04ec6e0c0:
    component is true;
  attribute fpga_dont_touch of bmg_72_e02664f04ec6e0c0:
    component is "true";
  attribute box_type of bmg_72_e02664f04ec6e0c0:
    component  is "black_box";
  component bmg_72_5ed93725c6f3d1db
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_5ed93725c6f3d1db:
    component is true;
  attribute fpga_dont_touch of bmg_72_5ed93725c6f3d1db:
    component is "true";
  attribute box_type of bmg_72_5ed93725c6f3d1db:
    component  is "black_box";
  component bmg_72_3d733db2a81768b0
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_3d733db2a81768b0:
    component is true;
  attribute fpga_dont_touch of bmg_72_3d733db2a81768b0:
    component is "true";
  attribute box_type of bmg_72_3d733db2a81768b0:
    component  is "black_box";
  component bmg_72_618ffcc3f0781f68
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_618ffcc3f0781f68:
    component is true;
  attribute fpga_dont_touch of bmg_72_618ffcc3f0781f68:
    component is "true";
  attribute box_type of bmg_72_618ffcc3f0781f68:
    component  is "black_box";
begin
  core_addr <= addr;
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_180432cd81ea5a8d")) generate
    core_instance0: bmg_72_180432cd81ea5a8d
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp1: if ((core_name0 = "bmg_72_8574240a262aac9a")) generate
    core_instance1: bmg_72_8574240a262aac9a
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp2: if ((core_name0 = "bmg_72_ce7e9961dfcc2802")) generate
    core_instance2: bmg_72_ce7e9961dfcc2802
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp3: if ((core_name0 = "bmg_72_e02664f04ec6e0c0")) generate
    core_instance3: bmg_72_e02664f04ec6e0c0
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp4: if ((core_name0 = "bmg_72_5ed93725c6f3d1db")) generate
    core_instance4: bmg_72_5ed93725c6f3d1db
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp5: if ((core_name0 = "bmg_72_3d733db2a81768b0")) generate
    core_instance5: bmg_72_3d733db2a81768b0
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp6: if ((core_name0 = "bmg_72_618ffcc3f0781f68")) generate
    core_instance6: bmg_72_618ffcc3f0781f68
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_1: if (latency <= 1) generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4670f4967f is
  port (
    d : in std_logic_vector((12 - 1) downto 0);
    q : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4670f4967f;


architecture behavior of delay_4670f4967f is
  signal d_1_22: std_logic_vector((12 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_08ed6107eb is
  port (
    in0 : in std_logic_vector((12 - 1) downto 0);
    in1 : in std_logic_vector((12 - 1) downto 0);
    in2 : in std_logic_vector((12 - 1) downto 0);
    in3 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((48 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_08ed6107eb;


architecture behavior of concat_08ed6107eb is
  signal in0_1_23: unsigned((12 - 1) downto 0);
  signal in1_1_27: unsigned((12 - 1) downto 0);
  signal in2_1_31: unsigned((12 - 1) downto 0);
  signal in3_1_35: unsigned((12 - 1) downto 0);
  signal y_2_1_concat: unsigned((48 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0c7cd7a34 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0c7cd7a34;


architecture behavior of concat_a0c7cd7a34 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_28d2c9d50c is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_28d2c9d50c;


architecture behavior of delay_28d2c9d50c is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (6 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(5);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e4b9fcaf02 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e4b9fcaf02;


architecture behavior of delay_e4b9fcaf02 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_a14e3dd1bd is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_a14e3dd1bd;


architecture behavior of delay_a14e3dd1bd is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_fca786f2ff is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((36 - 1) downto 0);
    d1 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_fca786f2ff;


architecture behavior of mux_fca786f2ff is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((36 - 1) downto 0);
  signal d1_1_27: std_logic_vector((36 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((36 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((36 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_5a12f8f9be is
  port (
    in0 : in std_logic_vector((19 - 1) downto 0);
    in1 : in std_logic_vector((19 - 1) downto 0);
    y : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_5a12f8f9be;


architecture behavior of concat_5a12f8f9be is
  signal in0_1_23: unsigned((19 - 1) downto 0);
  signal in1_1_27: unsigned((19 - 1) downto 0);
  signal y_2_1_concat: unsigned((38 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c615d93998 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c615d93998;


architecture behavior of concat_c615d93998 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((21 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_4a8cbc85ce is
  port (
    input_port : in std_logic_vector((20 - 1) downto 0);
    output_port : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_4a8cbc85ce;


architecture behavior of reinterpret_4a8cbc85ce is
  signal input_port_1_40: signed((20 - 1) downto 0);
  signal output_port_5_5_force: unsigned((20 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_d357e69fa3 is
  port (
    input_port : in std_logic_vector((21 - 1) downto 0);
    output_port : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_d357e69fa3;


architecture behavior of reinterpret_d357e69fa3 is
  signal input_port_1_40: unsigned((21 - 1) downto 0);
  signal output_port_5_5_force: signed((21 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_89dc141487 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_89dc141487;


architecture behavior of logical_89dc141487 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (2 - 1)) of std_logic;
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    '0',
    '0');
  signal latency_pipe_5_26_front_din: std_logic;
  signal latency_pipe_5_26_back: std_logic;
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal bit_2_27: std_logic;
  signal fully_2_1_bitnot: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(1);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          latency_pipe_5_26(i) <= latency_pipe_5_26(i-1);
        end loop;
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  bit_2_27 <= d0_1_24 and d1_1_27;
  fully_2_1_bitnot <= not bit_2_27;
  latency_pipe_5_26_front_din <= fully_2_1_bitnot;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= std_logic_to_vector(latency_pipe_5_26_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_f86ebb6084 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((20 - 1) downto 0);
    in2 : in std_logic_vector((20 - 1) downto 0);
    in3 : in std_logic_vector((20 - 1) downto 0);
    y : out std_logic_vector((80 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_f86ebb6084;


architecture behavior of concat_f86ebb6084 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((20 - 1) downto 0);
  signal in2_1_31: unsigned((20 - 1) downto 0);
  signal in3_1_35: unsigned((20 - 1) downto 0);
  signal y_2_1_concat: unsigned((80 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b366689086 is
  port (
    op : out std_logic_vector((19 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b366689086;


architecture behavior of constant_b366689086 is
begin
  op <= "0000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_b1e9d7c303 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_b1e9d7c303;


architecture behavior of logical_b1e9d7c303 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal bit_2_26: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bitnot: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  bit_2_26 <= d0_1_24 or d1_1_27;
  fully_2_1_bitnot <= not bit_2_26;
  y <= fully_2_1_bitnot;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_d930162434 is
  port (
    a : in std_logic_vector((4 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_d930162434;


architecture behavior of relational_d930162434 is
  signal a_1_31: unsigned((4 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_bd20dd351d is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_bd20dd351d;


architecture behavior of concat_bd20dd351d is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((2 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9a54e08c7c is
  port (
    input_port : in std_logic_vector((2 - 1) downto 0);
    output_port : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9a54e08c7c;


architecture behavior of reinterpret_9a54e08c7c is
  signal input_port_1_40: unsigned((2 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_713b6c5d29 is
  port (
    input_port : in std_logic_vector((20 - 1) downto 0);
    output_port : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_713b6c5d29;


architecture behavior of reinterpret_713b6c5d29 is
  signal input_port_1_40: unsigned((20 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_ce20fdf7b8 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((20 - 1) downto 0);
    d1 : in std_logic_vector((20 - 1) downto 0);
    y : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_ce20fdf7b8;


architecture behavior of mux_ce20fdf7b8 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((20 - 1) downto 0);
  signal d1_1_27: std_logic_vector((20 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((20 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "00000000000000000000",
    "00000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((20 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((20 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((20 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4822199898 is
  port (
    in0 : in std_logic_vector((38 - 1) downto 0);
    in1 : in std_logic_vector((38 - 1) downto 0);
    y : out std_logic_vector((76 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4822199898;


architecture behavior of concat_4822199898 is
  signal in0_1_23: unsigned((38 - 1) downto 0);
  signal in1_1_27: unsigned((38 - 1) downto 0);
  signal y_2_1_concat: unsigned((76 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4c449dd556 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4c449dd556;


architecture behavior of constant_4c449dd556 is
begin
  op <= "0000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_aab7b18c27 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_aab7b18c27;


architecture behavior of delay_aab7b18c27 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (6 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(5);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_d7d801964d is
  port (
    in0 : in std_logic_vector((12 - 1) downto 0);
    in1 : in std_logic_vector((12 - 1) downto 0);
    in2 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_d7d801964d;


architecture behavior of concat_d7d801964d is
  signal in0_1_23: unsigned((12 - 1) downto 0);
  signal in1_1_27: unsigned((12 - 1) downto 0);
  signal in2_1_31: unsigned((12 - 1) downto 0);
  signal y_2_1_concat: unsigned((36 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_87cc993d41 is
  port (
    d : in std_logic_vector((12 - 1) downto 0);
    q : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_87cc993d41;


architecture behavior of delay_87cc993d41 is
  signal d_1_22: std_logic_vector((12 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((12 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_452c4d3410 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_452c4d3410;


architecture behavior of concat_452c4d3410 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_1b04a69dde is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_1b04a69dde;


architecture behavior of delay_1b04a69dde is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (7 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(6);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 6 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_14a6a51cbc is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_14a6a51cbc;


architecture behavior of delay_14a6a51cbc is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (8 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(7);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 7 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_23d71a76f2 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_23d71a76f2;


architecture behavior of delay_23d71a76f2 is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4b00a70dea is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4b00a70dea;


architecture behavior of delay_4b00a70dea is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_6cd08a247e is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_6cd08a247e;


architecture behavior of counter_6cd08a247e is
  signal count_reg_20_23: unsigned((12 - 1) downto 0) := "000000000000";
begin
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if (ce = '1') then
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_0309b30f97 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_0309b30f97;


architecture behavior of logical_0309b30f97 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  type array_type_latency_pipe_5_26 is array (0 to (1 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    0 => "0");
  signal latency_pipe_5_26_front_din: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_back: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  latency_pipe_5_26_back <= latency_pipe_5_26(0);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  latency_pipe_5_26_front_din <= fully_2_1_bit;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= latency_pipe_5_26_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9e724c4b50 is
  port (
    in0 : in std_logic_vector((20 - 1) downto 0);
    in1 : in std_logic_vector((20 - 1) downto 0);
    y : out std_logic_vector((40 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9e724c4b50;


architecture behavior of concat_9e724c4b50 is
  signal in0_1_23: unsigned((20 - 1) downto 0);
  signal in1_1_27: unsigned((20 - 1) downto 0);
  signal y_2_1_concat: unsigned((40 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e6bc20c81b is
  port (
    in0 : in std_logic_vector((21 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((22 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e6bc20c81b;


architecture behavior of concat_e6bc20c81b is
  signal in0_1_23: unsigned((21 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((22 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_f0ca8483cb is
  port (
    input_port : in std_logic_vector((21 - 1) downto 0);
    output_port : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_f0ca8483cb;


architecture behavior of reinterpret_f0ca8483cb is
  signal input_port_1_40: signed((21 - 1) downto 0);
  signal output_port_5_5_force: unsigned((21 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_c84451c80b is
  port (
    input_port : in std_logic_vector((22 - 1) downto 0);
    output_port : out std_logic_vector((22 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_c84451c80b;


architecture behavior of reinterpret_c84451c80b is
  signal input_port_1_40: unsigned((22 - 1) downto 0);
  signal output_port_5_5_force: signed((22 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_fe87bb6ae4 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_fe87bb6ae4;


architecture behavior of logical_fe87bb6ae4 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (2 - 1)) of std_logic;
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    '0',
    '0');
  signal latency_pipe_5_26_front_din: std_logic;
  signal latency_pipe_5_26_back: std_logic;
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal bit_2_27: std_logic;
  signal fully_2_1_bitnot: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(1);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          latency_pipe_5_26(i) <= latency_pipe_5_26(i-1);
        end loop;
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  bit_2_27 <= d0_1_24 and d1_1_27 and d2_1_30;
  fully_2_1_bitnot <= not bit_2_27;
  latency_pipe_5_26_front_din <= fully_2_1_bitnot;
  latency_pipe_5_26_push_front_pop_back_en <= '1';
  y <= std_logic_to_vector(latency_pipe_5_26_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_356a264444 is
  port (
    in0 : in std_logic_vector((21 - 1) downto 0);
    in1 : in std_logic_vector((21 - 1) downto 0);
    in2 : in std_logic_vector((21 - 1) downto 0);
    in3 : in std_logic_vector((21 - 1) downto 0);
    y : out std_logic_vector((84 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_356a264444;


architecture behavior of concat_356a264444 is
  signal in0_1_23: unsigned((21 - 1) downto 0);
  signal in1_1_27: unsigned((21 - 1) downto 0);
  signal in2_1_31: unsigned((21 - 1) downto 0);
  signal in3_1_35: unsigned((21 - 1) downto 0);
  signal y_2_1_concat: unsigned((84 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity scale_97239b8ed2 is
  port (
    ip : in std_logic_vector((20 - 1) downto 0);
    op : out std_logic_vector((20 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end scale_97239b8ed2;


architecture behavior of scale_97239b8ed2 is
  signal ip_17_23: signed((20 - 1) downto 0);
begin
  ip_17_23 <= std_logic_vector_to_signed(ip);
  op <= signed_to_std_logic_vector(ip_17_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_299ca43e25 is
  port (
    input_port : in std_logic_vector((21 - 1) downto 0);
    output_port : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_299ca43e25;


architecture behavior of reinterpret_299ca43e25 is
  signal input_port_1_40: unsigned((21 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_46aae2a33a is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((21 - 1) downto 0);
    d1 : in std_logic_vector((21 - 1) downto 0);
    y : out std_logic_vector((21 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_46aae2a33a;


architecture behavior of mux_46aae2a33a is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((21 - 1) downto 0);
  signal d1_1_27: std_logic_vector((21 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((21 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000000000000",
    "000000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((21 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((21 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((21 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_83820b2faf is
  port (
    in0 : in std_logic_vector((37 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_83820b2faf;


architecture behavior of concat_83820b2faf is
  signal in0_1_23: unsigned((37 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((38 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_db4c53ade5 is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_db4c53ade5;


architecture behavior of reinterpret_db4c53ade5 is
  signal input_port_1_40: signed((37 - 1) downto 0);
  signal output_port_5_5_force: unsigned((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_2da6af93c2 is
  port (
    op : out std_logic_vector((35 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_2da6af93c2;


architecture behavior of constant_2da6af93c2 is
begin
  op <= "00000000000000000011111111111111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_620dd01637 is
  port (
    input_port : in std_logic_vector((38 - 1) downto 0);
    output_port : out std_logic_vector((38 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_620dd01637;


architecture behavior of reinterpret_620dd01637 is
  signal input_port_1_40: unsigned((38 - 1) downto 0);
  signal output_port_5_5_force: signed((38 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_ec14c62a89 is
  port (
    input_port : in std_logic_vector((35 - 1) downto 0);
    output_port : out std_logic_vector((35 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_ec14c62a89;


architecture behavior of reinterpret_ec14c62a89 is
  signal input_port_1_40: unsigned((35 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_5b4829fb41 is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_5b4829fb41;


architecture behavior of reinterpret_5b4829fb41 is
  signal input_port_1_40: unsigned((37 - 1) downto 0);
  signal output_port_5_5_force: signed((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_8e134646d3 is
  port (
    d : in std_logic_vector((37 - 1) downto 0);
    q : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_8e134646d3;


architecture behavior of delay_8e134646d3 is
  signal d_1_22: std_logic_vector((37 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_b28df1ab2e is
  port (
    in0 : in std_logic_vector((36 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_b28df1ab2e;


architecture behavior of concat_b28df1ab2e is
  signal in0_1_23: unsigned((36 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((36 - 1) downto 0);
  signal y_2_1_concat: unsigned((73 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_892b735f0d is
  port (
    input_port : in std_logic_vector((37 - 1) downto 0);
    output_port : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_892b735f0d;


architecture behavior of reinterpret_892b735f0d is
  signal input_port_1_40: unsigned((37 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_efdf1c3890 is
  port (
    input_port : in std_logic_vector((74 - 1) downto 0);
    output_port : out std_logic_vector((74 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_efdf1c3890;


architecture behavior of reinterpret_efdf1c3890 is
  signal input_port_1_40: unsigned((74 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c3ccc04d1a is
  port (
    in0 : in std_logic_vector((36 - 1) downto 0);
    in1 : in std_logic_vector((36 - 1) downto 0);
    y : out std_logic_vector((72 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c3ccc04d1a;


architecture behavior of concat_c3ccc04d1a is
  signal in0_1_23: unsigned((36 - 1) downto 0);
  signal in1_1_27: unsigned((36 - 1) downto 0);
  signal y_2_1_concat: unsigned((72 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_56d57d2c92 is
  port (
    in0 : in std_logic_vector((37 - 1) downto 0);
    in1 : in std_logic_vector((37 - 1) downto 0);
    y : out std_logic_vector((74 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_56d57d2c92;


architecture behavior of concat_56d57d2c92 is
  signal in0_1_23: unsigned((37 - 1) downto 0);
  signal in1_1_27: unsigned((37 - 1) downto 0);
  signal y_2_1_concat: unsigned((74 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mult_f295e5f0f2 is
  port (
    a : in std_logic_vector((18 - 1) downto 0);
    b : in std_logic_vector((18 - 1) downto 0);
    p : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mult_f295e5f0f2;


architecture behavior of mult_f295e5f0f2 is
  signal a_1_22: signed((18 - 1) downto 0);
  signal b_1_25: signed((18 - 1) downto 0);
  type array_type_op_mem_65_20 is array (0 to (2 - 1)) of signed((36 - 1) downto 0);
  signal op_mem_65_20: array_type_op_mem_65_20 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_65_20_front_din: signed((36 - 1) downto 0);
  signal op_mem_65_20_back: signed((36 - 1) downto 0);
  signal op_mem_65_20_push_front_pop_back_en: std_logic;
  signal mult_46_56: signed((36 - 1) downto 0);
begin
  a_1_22 <= std_logic_vector_to_signed(a);
  b_1_25 <= std_logic_vector_to_signed(b);
  op_mem_65_20_back <= op_mem_65_20(1);
  proc_op_mem_65_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_65_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_65_20(i) <= op_mem_65_20(i-1);
        end loop;
        op_mem_65_20(0) <= op_mem_65_20_front_din;
      end if;
    end if;
  end process proc_op_mem_65_20;
  mult_46_56 <= (a_1_22 * b_1_25);
  op_mem_65_20_front_din <= mult_46_56;
  op_mem_65_20_push_front_pop_back_en <= '1';
  p <= signed_to_std_logic_vector(op_mem_65_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_8dd4a43ef5 is
  port (
    a : in std_logic_vector((36 - 1) downto 0);
    b : in std_logic_vector((36 - 1) downto 0);
    s : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_8dd4a43ef5;


architecture behavior of addsub_8dd4a43ef5 is
  signal a_17_32: signed((36 - 1) downto 0);
  signal b_17_35: signed((36 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (2 - 1)) of signed((37 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_91_20_front_din: signed((37 - 1) downto 0);
  signal op_mem_91_20_back: signed((37 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (2 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_71_18: signed((37 - 1) downto 0);
  signal cast_71_22: signed((37 - 1) downto 0);
  signal internal_s_71_5_addsub: signed((37 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_signed(b);
  op_mem_91_20_back <= op_mem_91_20(1);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(1);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 1 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_71_18 <= s2s_cast(a_17_32, 34, 37, 34);
  cast_71_22 <= s2s_cast(b_17_35, 34, 37, 34);
  internal_s_71_5_addsub <= cast_71_18 - cast_71_22;
  op_mem_91_20_front_din <= internal_s_71_5_addsub;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_4ded11ba54 is
  port (
    a : in std_logic_vector((36 - 1) downto 0);
    b : in std_logic_vector((36 - 1) downto 0);
    s : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_4ded11ba54;


architecture behavior of addsub_4ded11ba54 is
  signal a_17_32: signed((36 - 1) downto 0);
  signal b_17_35: signed((36 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (2 - 1)) of signed((37 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_91_20_front_din: signed((37 - 1) downto 0);
  signal op_mem_91_20_back: signed((37 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (2 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    "0",
    "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: signed((37 - 1) downto 0);
  signal cast_69_22: signed((37 - 1) downto 0);
  signal internal_s_69_5_addsub: signed((37 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_signed(a);
  b_17_35 <= std_logic_vector_to_signed(b);
  op_mem_91_20_back <= op_mem_91_20(1);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_91_20(i) <= op_mem_91_20(i-1);
        end loop;
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(1);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        for i_x_000000 in 1 downto 1 loop 
          cout_mem_92_22(i_x_000000) <= cout_mem_92_22(i_x_000000-1);
        end loop;
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= s2s_cast(a_17_32, 34, 37, 34);
  cast_69_22 <= s2s_cast(b_17_35, 34, 37, 34);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  op_mem_91_20_front_din <= internal_s_69_5_addsub;
  op_mem_91_20_push_front_pop_back_en <= '1';
  cout_mem_92_22_front_din <= std_logic_vector_to_unsigned("0");
  cout_mem_92_22_push_front_pop_back_en <= '1';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= signed_to_std_logic_vector(op_mem_91_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_2d0f74b2c1 is
  port (
    d : in std_logic_vector((37 - 1) downto 0);
    q : out std_logic_vector((37 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_2d0f74b2c1;


architecture behavior of delay_2d0f74b2c1 is
  signal d_1_22: std_logic_vector((37 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000",
    "0000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((37 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9779a5cf83 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9779a5cf83;


architecture behavior of concat_9779a5cf83 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cda50df78a is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cda50df78a;


architecture behavior of constant_cda50df78a is
begin
  op <= "00";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity addsub_5e958c86e4 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    s : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end addsub_5e958c86e4;


architecture behavior of addsub_5e958c86e4 is
  signal a_17_32: unsigned((2 - 1) downto 0);
  signal b_17_35: unsigned((2 - 1) downto 0);
  type array_type_op_mem_91_20 is array (0 to (1 - 1)) of unsigned((2 - 1) downto 0);
  signal op_mem_91_20: array_type_op_mem_91_20 := (
    0 => "00");
  signal op_mem_91_20_front_din: unsigned((2 - 1) downto 0);
  signal op_mem_91_20_back: unsigned((2 - 1) downto 0);
  signal op_mem_91_20_push_front_pop_back_en: std_logic;
  type array_type_cout_mem_92_22 is array (0 to (1 - 1)) of unsigned((1 - 1) downto 0);
  signal cout_mem_92_22: array_type_cout_mem_92_22 := (
    0 => "0");
  signal cout_mem_92_22_front_din: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_back: unsigned((1 - 1) downto 0);
  signal cout_mem_92_22_push_front_pop_back_en: std_logic;
  signal prev_mode_93_22_next: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22: unsigned((3 - 1) downto 0);
  signal prev_mode_93_22_reg_i: std_logic_vector((3 - 1) downto 0);
  signal prev_mode_93_22_reg_o: std_logic_vector((3 - 1) downto 0);
  signal cast_69_18: unsigned((3 - 1) downto 0);
  signal cast_69_22: unsigned((3 - 1) downto 0);
  signal internal_s_69_5_addsub: unsigned((3 - 1) downto 0);
  signal cast_internal_s_83_3_convert: unsigned((2 - 1) downto 0);
begin
  a_17_32 <= std_logic_vector_to_unsigned(a);
  b_17_35 <= std_logic_vector_to_unsigned(b);
  op_mem_91_20_back <= op_mem_91_20(0);
  proc_op_mem_91_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_91_20_push_front_pop_back_en = '1')) then
        op_mem_91_20(0) <= op_mem_91_20_front_din;
      end if;
    end if;
  end process proc_op_mem_91_20;
  cout_mem_92_22_back <= cout_mem_92_22(0);
  proc_cout_mem_92_22: process (clk)
  is
    variable i_x_000000: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (cout_mem_92_22_push_front_pop_back_en = '1')) then
        cout_mem_92_22(0) <= cout_mem_92_22_front_din;
      end if;
    end if;
  end process proc_cout_mem_92_22;
  prev_mode_93_22_reg_i <= unsigned_to_std_logic_vector(prev_mode_93_22_next);
  prev_mode_93_22 <= std_logic_vector_to_unsigned(prev_mode_93_22_reg_o);
  prev_mode_93_22_reg_inst: entity work.synth_reg_w_init
    generic map (
      init_index => 2, 
      init_value => b"010", 
      latency => 1, 
      width => 3)
    port map (
      ce => ce, 
      clk => clk, 
      clr => clr, 
      i => prev_mode_93_22_reg_i, 
      o => prev_mode_93_22_reg_o);
  cast_69_18 <= u2u_cast(a_17_32, 0, 3, 0);
  cast_69_22 <= u2u_cast(b_17_35, 0, 3, 0);
  internal_s_69_5_addsub <= cast_69_18 + cast_69_22;
  cast_internal_s_83_3_convert <= u2u_cast(internal_s_69_5_addsub, 0, 2, 0);
  op_mem_91_20_push_front_pop_back_en <= '0';
  cout_mem_92_22_push_front_pop_back_en <= '0';
  prev_mode_93_22_next <= std_logic_vector_to_unsigned("000");
  s <= unsigned_to_std_logic_vector(cast_internal_s_83_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7eef56098d is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7eef56098d;


architecture behavior of concat_7eef56098d is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_09771002d6 is
  port (
    d : in std_logic_vector((9 - 1) downto 0);
    q : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_09771002d6;


architecture behavior of delay_09771002d6 is
  signal d_1_22: std_logic_vector((9 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000");
  signal op_mem_20_24_front_din: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_pipeline is
    generic (
        old_width   : integer := 16;
        old_bin_pt  : integer := 4;
        old_arith   : integer := xlUnsigned;
        new_width   : integer := 8;
        new_bin_pt  : integer := 2;
        new_arith   : integer := xlUnsigned;
        en_width    : integer := 1;
        en_bin_pt   : integer := 0;
        en_arith    : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow    : integer := xlWrap;
        latency     : integer := 1);
    port (
        din : in std_logic_vector (old_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        result : out std_logic_vector (new_width-1 downto 0));
end convert_pipeline;
architecture behavior of convert_pipeline is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i           : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    constant fp_width : integer := old_width + 2;
    constant fp_bin_pt : integer := old_bin_pt;
    constant fp_arith : integer := old_arith;
    constant q_width : integer := (old_width + 2) + (new_bin_pt - old_bin_pt);
    constant q_bin_pt : integer := new_bin_pt;
    constant q_arith : integer := old_arith;
    signal full_precision_result_in, full_precision_result_out
        : std_logic_vector(fp_width-1 downto 0);
    signal quantized_result_in, quantized_result_out
        : std_logic_vector(q_width-1 downto 0);
    signal result_in : std_logic_vector(new_width-1 downto 0):= (others => '0');
    signal internal_ce : std_logic;
begin
    internal_ce <= ce and en(0);

    fp_result : process (din)
    begin
        full_precision_result_in <= cast(din, old_bin_pt,
                                         fp_width, fp_bin_pt, fp_arith);
    end process;
    latency_fpr : if (latency > 2)
    generate
        reg_fpr : synth_reg
            generic map ( width => fp_width,
                          latency => 1)
            port map (i => full_precision_result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => full_precision_result_out);
    end generate;
    no_latency_fpr : if (latency < 3)
    generate
        full_precision_result_out <= full_precision_result_in;
    end generate;
    xlround_generate : if (quantization = xlRound)
    generate
      xlround_result : process (full_precision_result_out)
      begin
          quantized_result_in <= round_towards_inf(full_precision_result_out,
                                                   fp_width, fp_bin_pt,
                                                   fp_arith, q_width, q_bin_pt,
                                                   q_arith);
      end process;
    end generate;
    xlroundbanker_generate : if (quantization = xlRoundBanker)
    generate
      xlroundbanker_result : process (full_precision_result_out)
      begin
          quantized_result_in <= round_towards_even(full_precision_result_out,
                                                   fp_width, fp_bin_pt,
                                                   fp_arith, q_width, q_bin_pt,
                                                   q_arith);
      end process;
    end generate;
    xltruncate_generate : if (quantization = xlTruncate)
    generate
      xltruncate_result : process (full_precision_result_out)
      begin
          quantized_result_in <= trunc(full_precision_result_out,
                                       fp_width, fp_bin_pt,
                                       fp_arith, q_width, q_bin_pt,
                                       q_arith);
      end process;
    end generate;
    latency_qr : if (latency > 1)
    generate
        reg_qr : synth_reg
            generic map ( width => q_width,
                          latency => 1)
            port map (i => quantized_result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => quantized_result_out);
    end generate;
    no_latency_qr : if (latency < 2)
    generate
        quantized_result_out <= quantized_result_in;
    end generate;
    xlsaturate_generate : if (overflow = xlSaturate)
    generate
      xlsaturate_result : process (quantized_result_out)
      begin
          result_in <= saturation_arith(quantized_result_out, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
      end process;
    end generate;
    xlwrap_generate : if (overflow = xlWrap)
    generate
      xlwrap_result : process (quantized_result_out)
      begin
          result_in <= wrap_arith(quantized_result_out, q_width, q_bin_pt,
                                  q_arith, new_width, new_bin_pt, new_arith);
      end process;
    end generate;
    latency_gt_3 : if (latency > 3)
    generate
        reg_out : synth_reg
            generic map ( width => new_width,
                          latency => latency-2)
            port map (i => result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => result);
    end generate;
    latency_lt_4 : if ((latency < 4) and (latency > 0))
    generate
        reg_out : synth_reg
            generic map ( width => new_width,
                          latency => 1)
            port map (i => result_in,
                      ce => internal_ce,
                      clr => clr,
                      clk => clk,
                      o => result);
    end generate;
    latency0 : if (latency = 0)
    generate
        result <= result_in;
    end generate latency0;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert_pipeline is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din  : in std_logic_vector (din_width-1 downto 0);
        en   : in std_logic_vector (en_width-1 downto 0);
        ce   : in std_logic;
        clr  : in std_logic;
        clk  : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert_pipeline;
architecture behavior of xlconvert_pipeline is
    component convert_pipeline
        generic (
            old_width    : integer := 16;
            old_bin_pt   : integer := 4;
            old_arith    : integer := xlUnsigned;
            new_width    : integer := 8;
            new_bin_pt   : integer := 2;
            new_arith    : integer := xlUnsigned;
            en_width     : integer := 1;
            en_bin_pt    : integer := 0;
            en_arith     : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap;
            latency      : integer := 1);
        port (
            din    : in std_logic_vector (din_width-1 downto 0);
            en     : in std_logic_vector (en_width-1 downto 0);
            ce     : in std_logic;
            clr    : in std_logic;
            clk    : in std_logic;
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
   begin
      convert : convert_pipeline
        generic map (
          old_width   => din_width,
          old_bin_pt  => din_bin_pt,
          old_arith   => din_arith,
          new_width   => dout_width,
          new_bin_pt  => dout_bin_pt,
          new_arith   => dout_arith,
          en_width    => en_width,
          en_bin_pt   => en_bin_pt,
          en_arith    => en_arith,
          quantization => quantization,
          overflow    => overflow,
          latency     => latency)
        port map (
          din => din,
          en => en,
          ce => ce,
          clr => clr,
          clk => clk,
          result => dout);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_6104cbef7a is
  port (
    d : in std_logic_vector((9 - 1) downto 0);
    q : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_6104cbef7a;


architecture behavior of delay_6104cbef7a is
  signal d_1_22: std_logic_vector((9 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000",
    "000000000");
  signal op_mem_20_24_front_din: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((9 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_3ffe3e5660 is
  port (
    d : in std_logic_vector((73 - 1) downto 0);
    q : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_3ffe3e5660;


architecture behavior of delay_3ffe3e5660 is
  signal d_1_22: std_logic_vector((73 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_b6092ad150 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_b6092ad150;


architecture behavior of delay_b6092ad150 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_206b7f76d8 is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_206b7f76d8;


architecture behavior of negate_206b7f76d8 is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (1 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    0 => "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(0);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  internal_ip_40_3_convert <= std_logic_vector_to_signed(convert_type(signed_to_std_logic_vector(internal_ip_join_30_1), 19, 17, xlSigned, 18, 17, xlSigned, xlTruncate, xlSaturate));
  op_mem_48_20_front_din <= internal_ip_40_3_convert;
  op_mem_48_20_push_front_pop_back_en <= '1';
  op <= signed_to_std_logic_vector(op_mem_48_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_1896e7760c is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_1896e7760c;


architecture behavior of mux_1896e7760c is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000000000",
    "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4e7d828d94 is
  port (
    d : in std_logic_vector((73 - 1) downto 0);
    q : out std_logic_vector((73 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4e7d828d94;


architecture behavior of delay_4e7d828d94 is
  signal d_1_22: std_logic_vector((73 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000",
    "0000000000000000000000000000000000000000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((73 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlpassthrough is
    generic (
        din_width    : integer := 16;
        dout_width   : integer := 16
        );
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlpassthrough;
architecture passthrough_arch of xlpassthrough is
begin
  dout <= din;
end passthrough_arch;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_8f386731a6 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_8f386731a6;


architecture behavior of counter_8f386731a6 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((12 - 1) downto 0) := "000000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((13 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_cfdc93535e is
  port (
    in0 : in std_logic_vector((40 - 1) downto 0);
    in1 : in std_logic_vector((40 - 1) downto 0);
    y : out std_logic_vector((80 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_cfdc93535e;


architecture behavior of concat_cfdc93535e is
  signal in0_1_23: unsigned((40 - 1) downto 0);
  signal in1_1_27: unsigned((40 - 1) downto 0);
  signal y_2_1_concat: unsigned((80 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_faa52967c8 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_faa52967c8;


architecture behavior of delay_faa52967c8 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (8 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(7);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 7 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_67ad97ca70 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_67ad97ca70;


architecture behavior of constant_67ad97ca70 is
begin
  op <= "0001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_145086465d is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_145086465d;


architecture behavior of constant_145086465d is
begin
  op <= "1000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_230536be32 is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((4 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_230536be32;


architecture behavior of counter_230536be32 is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((4 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((4 - 1) downto 0);
  signal count_reg_20_23: unsigned((4 - 1) downto 0) := "0000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((6 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((6 - 1) downto 0);
  signal count_reg_join_48_3: signed((6 - 1) downto 0);
  signal count_reg_join_44_1: signed((6 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((4 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 6, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 6, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 4, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_4d3cfceaf4 is
  port (
    a : in std_logic_vector((4 - 1) downto 0);
    b : in std_logic_vector((4 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_4d3cfceaf4;


architecture behavior of relational_4d3cfceaf4 is
  signal a_1_31: unsigned((4 - 1) downto 0);
  signal b_1_34: unsigned((4 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0c0a0420a6 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0c0a0420a6;


architecture behavior of delay_0c0a0420a6 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0341f7be44 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0341f7be44;


architecture behavior of delay_0341f7be44 is
  signal d_1_22: std_logic;
begin
  d_1_22 <= d(0);
  q <= std_logic_to_vector(d_1_22);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_6068817c97 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_6068817c97;


architecture behavior of counter_6068817c97 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((4 - 1) downto 0) := "0000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((5 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("0001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e774b32dc9 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e774b32dc9;


architecture behavior of concat_e774b32dc9 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_811dd91a3d is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((10 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_811dd91a3d;


architecture behavior of concat_811dd91a3d is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((10 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4fd36a24a3 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4fd36a24a3;


architecture behavior of concat_4fd36a24a3 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_cf4f99539f is
  port (
    d : in std_logic_vector((10 - 1) downto 0);
    q : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_cf4f99539f;


architecture behavior of delay_cf4f99539f is
  signal d_1_22: std_logic_vector((10 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000000000");
  signal op_mem_20_24_front_din: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_325391d82e is
  port (
    d : in std_logic_vector((10 - 1) downto 0);
    q : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_325391d82e;


architecture behavior of delay_325391d82e is
  signal d_1_22: std_logic_vector((10 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000000",
    "0000000000");
  signal op_mem_20_24_front_din: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((10 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a7e2bb9e12 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a7e2bb9e12;


architecture behavior of constant_a7e2bb9e12 is
begin
  op <= "01";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xldpram_fft_astro_devel_core is
  generic (
    core_name0: string := "";
    c_width_a: integer := 13;
    c_address_width_a: integer := 4;
    c_width_b: integer := 13;
    c_address_width_b: integer := 4;
    c_has_sinita: integer := 0;
    c_has_sinitb: integer := 0;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width_a - 1 downto 0);
    addra: in std_logic_vector(c_address_width_a - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    a_ce: in std_logic;
    a_clk: in std_logic;
    rsta: in std_logic_vector(0 downto 0) := (others => '0');
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    douta: out std_logic_vector(c_width_a - 1 downto 0);
    dinb: in std_logic_vector(c_width_b - 1 downto 0);
    addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
    web: in std_logic_vector(0 downto 0);
    b_ce: in std_logic;
    b_clk: in std_logic;
    rstb: in std_logic_vector(0 downto 0) := (others => '0');
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    doutb: out std_logic_vector(c_width_b - 1 downto 0)
  );
end xldpram_fft_astro_devel_core;
architecture behavior of xldpram_fft_astro_devel_core is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;

  signal core_addra: std_logic_vector(c_address_width_a - 1 downto 0);
  signal core_addrb: std_logic_vector(c_address_width_b - 1 downto 0);
  signal core_dina, core_douta, dly_douta:
    std_logic_vector(c_width_a - 1 downto 0);
  signal core_dinb, core_doutb, dly_doutb:
    std_logic_vector(c_width_b - 1 downto 0);
  signal core_wea, core_web: std_logic;
  signal core_a_ce, core_b_ce: std_logic;
  signal sinita, sinitb: std_logic;

  component bmg_72_9f585cf1e3329833
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_9f585cf1e3329833:
    component is true;
  attribute fpga_dont_touch of bmg_72_9f585cf1e3329833:
    component is "true";
  attribute box_type of bmg_72_9f585cf1e3329833:
    component  is "black_box";
  component bmg_72_15a84ff1ccdd3419
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_15a84ff1ccdd3419:
    component is true;
  attribute fpga_dont_touch of bmg_72_15a84ff1ccdd3419:
    component is "true";
  attribute box_type of bmg_72_15a84ff1ccdd3419:
    component  is "black_box";
  component bmg_72_9d950569c0d7f9e8
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_9d950569c0d7f9e8:
    component is true;
  attribute fpga_dont_touch of bmg_72_9d950569c0d7f9e8:
    component is "true";
  attribute box_type of bmg_72_9d950569c0d7f9e8:
    component  is "black_box";
begin
  core_addra <= addra;
  core_dina <= dina;
  douta <= dly_douta;
  core_wea <= wea(0);
  core_a_ce <= a_ce and ena(0);
  sinita <= rsta(0) and a_ce;

  core_addrb <= addrb;
  core_dinb <= dinb;
  doutb <= dly_doutb;
  core_web <= web(0);
  core_b_ce <= b_ce and enb(0);
  sinitb <= rstb(0) and b_ce;
  comp0: if ((core_name0 = "bmg_72_9f585cf1e3329833")) generate
    core_instance0: bmg_72_9f585cf1e3329833
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_15a84ff1ccdd3419")) generate
    core_instance1: bmg_72_15a84ff1ccdd3419
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp2: if ((core_name0 = "bmg_72_9d950569c0d7f9e8")) generate
    core_instance2: bmg_72_9d950569c0d7f9e8
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  latency_test: if (latency > 2) generate
    regA: synth_reg
      generic map (
        width => c_width_a,
        latency => latency - 2
      )
      port map (
        i => core_douta,
        ce => core_a_ce,
        clr => '0',
        clk => a_clk,
        o => dly_douta
      );
    regB: synth_reg
      generic map (
        width => c_width_b,
        latency => latency - 2
      )
      port map (
        i => core_doutb,
        ce => core_b_ce,
        clr => '0',
        clk => b_clk,
        o => dly_doutb
      );
  end generate;
  latency1: if (latency <= 2) generate
    dly_douta <= core_douta;
    dly_doutb <= core_doutb;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_95b0f967bc is
  port (
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_95b0f967bc;


architecture behavior of constant_95b0f967bc is
begin
  op <= "000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a1c496ea88 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a1c496ea88;


architecture behavior of constant_a1c496ea88 is
begin
  op <= "001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_822933f89b is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_822933f89b;


architecture behavior of constant_822933f89b is
begin
  op <= "000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_469094441c is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_469094441c;


architecture behavior of constant_469094441c is
begin
  op <= "100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_ed7367cb5c is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((3 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_ed7367cb5c;


architecture behavior of counter_ed7367cb5c is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((3 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((3 - 1) downto 0);
  signal count_reg_20_23: unsigned((3 - 1) downto 0) := "000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((5 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((5 - 1) downto 0);
  signal count_reg_join_48_3: signed((5 - 1) downto 0);
  signal count_reg_join_44_1: signed((5 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((3 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 5, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("00001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 5, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 3, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_8fc7f5539b is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_8fc7f5539b;


architecture behavior of relational_8fc7f5539b is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_47b317dab6 is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_47b317dab6;


architecture behavior of relational_47b317dab6 is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_191d4874ab is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_191d4874ab;


architecture behavior of counter_191d4874ab is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((3 - 1) downto 0) := "000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((4 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0fa71d0d3 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    in10 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0fa71d0d3;


architecture behavior of concat_a0fa71d0d3 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal in10_1_63: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((11 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  in10_1_63 <= std_logic_vector_to_unsigned(in10);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59) & unsigned_to_std_logic_vector(in10_1_63));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9769d05421 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((11 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9769d05421;


architecture behavior of concat_9769d05421 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((11 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7ad1e33701 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((10 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7ad1e33701;


architecture behavior of concat_7ad1e33701 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((10 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0604807f72 is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0604807f72;


architecture behavior of constant_0604807f72 is
begin
  op <= "10000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_046d743d02 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((10 - 1) downto 0);
    d1 : in std_logic_vector((11 - 1) downto 0);
    y : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_046d743d02;


architecture behavior of mux_046d743d02 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((10 - 1) downto 0);
  signal d1_1_27: std_logic_vector((11 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((11 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "00000000000",
    "00000000000");
  signal pipe_16_22_front_din: std_logic_vector((11 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((11 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((11 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 11, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8ddc079e9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8ddc079e9;


architecture behavior of constant_e8ddc079e9 is
begin
  op <= "10";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_38898c80c0 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_38898c80c0;


architecture behavior of delay_38898c80c0 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_e095645f0c is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((2 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_e095645f0c;


architecture behavior of counter_e095645f0c is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((2 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((2 - 1) downto 0);
  signal count_reg_20_23: unsigned((2 - 1) downto 0) := "00";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((4 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((4 - 1) downto 0);
  signal count_reg_join_48_3: signed((4 - 1) downto 0);
  signal count_reg_join_44_1: signed((4 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((2 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 4, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("0001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 4, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 2, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5f1eb17108 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5f1eb17108;


architecture behavior of relational_5f1eb17108 is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_f9928864ea is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_f9928864ea;


architecture behavior of relational_f9928864ea is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_363af54ff2 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_363af54ff2;


architecture behavior of counter_363af54ff2 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((2 - 1) downto 0) := "00";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((3 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "00";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("01");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ef66525e56 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    in8 : in std_logic_vector((1 - 1) downto 0);
    in9 : in std_logic_vector((1 - 1) downto 0);
    in10 : in std_logic_vector((1 - 1) downto 0);
    in11 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ef66525e56;


architecture behavior of concat_ef66525e56 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal in8_1_55: unsigned((1 - 1) downto 0);
  signal in9_1_59: unsigned((1 - 1) downto 0);
  signal in10_1_63: unsigned((1 - 1) downto 0);
  signal in11_1_68: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((12 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  in8_1_55 <= std_logic_vector_to_unsigned(in8);
  in9_1_59 <= std_logic_vector_to_unsigned(in9);
  in10_1_63 <= std_logic_vector_to_unsigned(in10);
  in11_1_68 <= std_logic_vector_to_unsigned(in11);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51) & unsigned_to_std_logic_vector(in8_1_55) & unsigned_to_std_logic_vector(in9_1_59) & unsigned_to_std_logic_vector(in10_1_63) & unsigned_to_std_logic_vector(in11_1_68));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_118109a960 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_118109a960;


architecture behavior of concat_118109a960 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((12 - 1) downto 0);
  signal y_2_1_concat: unsigned((13 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_8503582fb5 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((11 - 1) downto 0);
    y : out std_logic_vector((13 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_8503582fb5;


architecture behavior of concat_8503582fb5 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((11 - 1) downto 0);
  signal y_2_1_concat: unsigned((13 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_49cb1051e0 is
  port (
    d : in std_logic_vector((11 - 1) downto 0);
    q : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_49cb1051e0;


architecture behavior of delay_49cb1051e0 is
  signal d_1_22: std_logic_vector((11 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000000000");
  signal op_mem_20_24_front_din: std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((11 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e054d850c5 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e054d850c5;


architecture behavior of constant_e054d850c5 is
begin
  op <= "100000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_efb9621913 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((11 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_efb9621913;


architecture behavior of mux_efb9621913 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((11 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (2 - 1)) of std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000",
    "000000000000");
  signal pipe_16_22_front_din: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((12 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(1);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 12, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_223a0f3237 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_223a0f3237;


architecture behavior of counter_223a0f3237 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((1 - 1) downto 0) := "0";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((2 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("1");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity negate_155cd8ddf7 is
  port (
    ip : in std_logic_vector((18 - 1) downto 0);
    op : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end negate_155cd8ddf7;


architecture behavior of negate_155cd8ddf7 is
  signal ip_18_25: signed((18 - 1) downto 0);
  type array_type_op_mem_48_20 is array (0 to (3 - 1)) of signed((18 - 1) downto 0);
  signal op_mem_48_20: array_type_op_mem_48_20 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_48_20_front_din: signed((18 - 1) downto 0);
  signal op_mem_48_20_back: signed((18 - 1) downto 0);
  signal op_mem_48_20_push_front_pop_back_en: std_logic;
  signal cast_35_24: signed((19 - 1) downto 0);
  signal internal_ip_35_9_neg: signed((19 - 1) downto 0);
  signal internal_ip_join_30_1: signed((19 - 1) downto 0);
  signal internal_ip_40_3_convert: signed((18 - 1) downto 0);
begin
  ip_18_25 <= std_logic_vector_to_signed(ip);
  op_mem_48_20_back <= op_mem_48_20(2);
  proc_op_mem_48_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_48_20_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_48_20(i) <= op_mem_48_20(i-1);
        end loop;
        op_mem_48_20(0) <= op_mem_48_20_front_din;
      end if;
    end if;
  end process proc_op_mem_48_20;
  cast_35_24 <= s2s_cast(ip_18_25, 17, 19, 17);
  internal_ip_35_9_neg <=  -cast_35_24;
  proc_if_30_1: process (internal_ip_35_9_neg)
  is
  begin
    if false then
      internal_ip_join_30_1 <= std_logic_vector_to_signed("0000000000000000000");
    else 
      internal_ip_join_30_1 <= internal_ip_35_9_neg;
    end if;
  end process proc_if_30_1;
  internal_ip_40_3_convert <= std_logic_vector_to_signed(convert_type(signed_to_std_logic_vector(internal_ip_join_30_1), 19, 17, xlSigned, 18, 17, xlSigned, xlTruncate, xlSaturate));
  op_mem_48_20_front_din <= internal_ip_40_3_convert;
  op_mem_48_20_push_front_pop_back_en <= '1';
  op <= signed_to_std_logic_vector(op_mem_48_20_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_328e8ebbb5 is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_328e8ebbb5;


architecture behavior of delay_328e8ebbb5 is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (3 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(2);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 2 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_dbbe492743 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_dbbe492743;


architecture behavior of delay_dbbe492743 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (9 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(8);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 8 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_621a1c5abf is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_621a1c5abf;


architecture behavior of mux_621a1c5abf is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (6 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(5);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        for i in 5 downto 1 loop 
          pipe_16_22(i) <= pipe_16_22(i-1);
        end loop;
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_43bd805056 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_43bd805056;


architecture behavior of delay_43bd805056 is
  signal d_1_22: std_logic_vector((1 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0",
    "0",
    "0",
    "0",
    "0");
  signal op_mem_20_24_front_din: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((1 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_c462a80bee is
  port (
    d : in std_logic_vector((18 - 1) downto 0);
    q : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_c462a80bee;


architecture behavior of delay_c462a80bee is
  signal d_1_22: std_logic_vector((18 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000",
    "000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((18 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_181e58d842 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((18 - 1) downto 0);
    d1 : in std_logic_vector((18 - 1) downto 0);
    y : out std_logic_vector((18 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_181e58d842;


architecture behavior of mux_181e58d842 is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((18 - 1) downto 0);
  signal d1_1_27: std_logic_vector((18 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "000000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((18 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal unregy_join_6_1: std_logic_vector((18 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_6b1adb5d55 is
  port (
    input_port : in std_logic_vector((11 - 1) downto 0);
    output_port : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_6b1adb5d55;


architecture behavior of reinterpret_6b1adb5d55 is
  signal input_port_1_40: unsigned((11 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_b754317574 is
  port (
    input_port : in std_logic_vector((9 - 1) downto 0);
    output_port : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_b754317574;


architecture behavior of reinterpret_b754317574 is
  signal input_port_1_40: unsigned((9 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_88cfa744f5 is
  port (
    in0 : in std_logic_vector((9 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    in2 : in std_logic_vector((9 - 1) downto 0);
    in3 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_88cfa744f5;


architecture behavior of concat_88cfa744f5 is
  signal in0_1_23: unsigned((9 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal in2_1_31: unsigned((9 - 1) downto 0);
  signal in3_1_35: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((36 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7c91b1b314 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7c91b1b314;


architecture behavior of constant_7c91b1b314 is
begin
  op <= "000000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd28b32bf8 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd28b32bf8;


architecture behavior of constant_fd28b32bf8 is
begin
  op <= "000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_a0220fdf9f is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((12 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_a0220fdf9f;


architecture behavior of counter_a0220fdf9f is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((12 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((12 - 1) downto 0);
  signal count_reg_20_23: unsigned((12 - 1) downto 0) := "000000000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((14 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((14 - 1) downto 0);
  signal count_reg_join_48_3: signed((14 - 1) downto 0);
  signal count_reg_join_44_1: signed((14 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((12 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 14, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("00000000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 14, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 12, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_d36fe12c1c is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_d36fe12c1c;


architecture behavior of relational_d36fe12c1c is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_acb3c05dd0 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_acb3c05dd0;


architecture behavior of relational_acb3c05dd0 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e18fb31a3d is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e18fb31a3d;


architecture behavior of delay_e18fb31a3d is
  signal d_1_22: std_logic;
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic;
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    '0',
    '0');
  signal op_mem_20_24_front_din: std_logic;
  signal op_mem_20_24_back: std_logic;
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d(0);
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= std_logic_to_vector(op_mem_20_24_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_7439478232 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_7439478232;


architecture behavior of delay_7439478232 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (5 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(4);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 4 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_e4b8f9ed4e is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_e4b8f9ed4e;


architecture behavior of counter_e4b8f9ed4e is
  signal count_reg_20_23: unsigned((11 - 1) downto 0) := "00000000000";
begin
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if (ce = '1') then
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("00000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e6f5ee726b is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e6f5ee726b;


architecture behavior of concat_e6f5ee726b is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((2 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_4a9a9a25a3 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_4a9a9a25a3;


architecture behavior of concat_4a9a9a25a3 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((2 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_6160d7387c is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_6160d7387c;


architecture behavior of concat_6160d7387c is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((3 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4ce33ca7e7 is
  port (
    d : in std_logic_vector((2 - 1) downto 0);
    q : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4ce33ca7e7;


architecture behavior of delay_4ce33ca7e7 is
  signal d_1_22: std_logic_vector((2 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00");
  signal op_mem_20_24_front_din: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_fcebea29b9 is
  port (
    d : in std_logic_vector((2 - 1) downto 0);
    q : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_fcebea29b9;


architecture behavior of delay_fcebea29b9 is
  signal d_1_22: std_logic_vector((2 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "00",
    "00");
  signal op_mem_20_24_front_din: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((2 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.6 VHDL source file.
--
-- Copyright(C) 2013 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2013 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldpram_dist_fft_astro_devel_core is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    addr_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width - 1 downto 0);
    addra: in std_logic_vector(addr_width - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    a_ce: in std_logic;
    a_clk: in std_logic;
    douta: out std_logic_vector(c_width - 1 downto 0);
    addrb: in std_logic_vector(addr_width - 1 downto 0);
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    b_ce: in std_logic;
    b_clk: in std_logic;
    doutb: out std_logic_vector(c_width - 1 downto 0)
  );
end xldpram_dist_fft_astro_devel_core ;
architecture behavior of xldpram_dist_fft_astro_devel_core is
  component synth_reg is
    generic (
      width: integer := 8;
      latency: integer := 1
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  constant num_extra_addr_bits: integer := (c_address_width - addr_width);
  signal core_addra, core_addrb: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_in, core_douta, core_doutb: std_logic_vector(c_width - 1 downto 0);
  signal reg_douta, reg_doutb: std_logic_vector(c_width - 1 downto 0);
  signal core_we: std_logic_vector(0 downto 0);
  signal core_cea, core_ceb: std_logic;
  component dmg_72_505931c5b3ea228e
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_505931c5b3ea228e:
    component is true;
  attribute fpga_dont_touch of dmg_72_505931c5b3ea228e:
    component is "true";
  attribute box_type of dmg_72_505931c5b3ea228e:
    component  is "black_box";
  component dmg_72_d20b02a9f8239c7a
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_d20b02a9f8239c7a:
    component is true;
  attribute fpga_dont_touch of dmg_72_d20b02a9f8239c7a:
    component is "true";
  attribute box_type of dmg_72_d20b02a9f8239c7a:
    component  is "black_box";
  component dmg_72_efdf1b1b05926829
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_efdf1b1b05926829:
    component is true;
  attribute fpga_dont_touch of dmg_72_efdf1b1b05926829:
    component is "true";
  attribute box_type of dmg_72_efdf1b1b05926829:
    component  is "black_box";
  component dmg_72_1c323e86177437db
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      d: in std_logic_vector(c_width - 1 downto 0);
      we: in std_logic;
      dpra: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0);
      dpo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_1c323e86177437db:
    component is true;
  attribute fpga_dont_touch of dmg_72_1c323e86177437db:
    component is "true";
  attribute box_type of dmg_72_1c323e86177437db:
    component  is "black_box";
begin
  need_to_pad_addr : if num_extra_addr_bits > 0 generate
      core_addra(c_address_width - 1 downto addr_width) <= (others => '0');
      core_addra(addr_width - 1 downto 0) <= addra;
      core_addrb(c_address_width - 1 downto addr_width) <= (others => '0');
      core_addrb(addr_width - 1 downto 0) <= addrb;
  end generate;
  no_need_to_pad_addr: if num_extra_addr_bits = 0 generate
    core_addra <= addra;
    core_addrb <= addrb;
  end generate;
  douta <= reg_douta;
  doutb <= reg_doutb;
  core_cea <= a_ce and ena(0);
  core_ceb <= b_ce and enb(0);
  core_we(0) <= wea(0) and core_cea;
  registered_dpram : if latency > 0 generate
    output_rega: synth_reg
      generic map (
        width   => c_width,
        latency => latency
      )
      port map (
        i   => core_douta,
        ce  => core_cea,
        clr => '0',
        clk => a_clk,
        o   => reg_douta
      );
    output_regb: synth_reg
      generic map (
        width   => c_width,
        latency => latency
      )
      port map (
        i   => core_doutb,
        ce  => core_ceb,
        clr => '0',
        clk => b_clk,
        o   => reg_doutb
      );
  end generate;
  nonregistered_ram : if latency = 0 generate
    reg_douta <= core_douta;
    reg_doutb <= core_doutb;
  end generate;
  comp0: if ((core_name0 = "dmg_72_505931c5b3ea228e")) generate
    core_instance0: dmg_72_505931c5b3ea228e
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "dmg_72_d20b02a9f8239c7a")) generate
    core_instance1: dmg_72_d20b02a9f8239c7a
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp2: if ((core_name0 = "dmg_72_efdf1b1b05926829")) generate
    core_instance2: dmg_72_efdf1b1b05926829
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
  comp3: if ((core_name0 = "dmg_72_1c323e86177437db")) generate
    core_instance3: dmg_72_1c323e86177437db
      port map (
        a => core_addra,
        clk => a_clk,
        d => dina,
        we => core_we(0),
        dpra => core_addrb,
        spo => core_douta,
        dpo => core_doutb
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_e262000247 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_e262000247;


architecture behavior of delay_e262000247 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1024 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1023);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1023 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_118598964d is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_118598964d;


architecture behavior of constant_118598964d is
begin
  op <= "00000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a3923dd146 is
  port (
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a3923dd146;


architecture behavior of constant_a3923dd146 is
begin
  op <= "00000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_b5e433c475 is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((11 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_b5e433c475;


architecture behavior of counter_b5e433c475 is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((11 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((11 - 1) downto 0);
  signal count_reg_20_23: unsigned((11 - 1) downto 0) := "00000000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((13 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((13 - 1) downto 0);
  signal count_reg_join_48_3: signed((13 - 1) downto 0);
  signal count_reg_join_44_1: signed((13 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((11 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 13, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("0000000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 13, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 11, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_2147430058 is
  port (
    a : in std_logic_vector((11 - 1) downto 0);
    b : in std_logic_vector((11 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_2147430058;


architecture behavior of relational_2147430058 is
  signal a_1_31: unsigned((11 - 1) downto 0);
  signal b_1_34: unsigned((11 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_b4b277ae0f is
  port (
    a : in std_logic_vector((11 - 1) downto 0);
    b : in std_logic_vector((11 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_b4b277ae0f;


architecture behavior of relational_b4b277ae0f is
  signal a_1_31: unsigned((11 - 1) downto 0);
  signal b_1_34: unsigned((11 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_21896c7599 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((11 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_21896c7599;


architecture behavior of counter_21896c7599 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((11 - 1) downto 0) := "00000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((12 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "00000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("00000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_949f038a6d is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_949f038a6d;


architecture behavior of concat_949f038a6d is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_54d5af2115 is
  port (
    d : in std_logic_vector((3 - 1) downto 0);
    q : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_54d5af2115;


architecture behavior of delay_54d5af2115 is
  signal d_1_22: std_logic_vector((3 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000");
  signal op_mem_20_24_front_din: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_6edcd04662 is
  port (
    d : in std_logic_vector((3 - 1) downto 0);
    q : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_6edcd04662;


architecture behavior of delay_6edcd04662 is
  signal d_1_22: std_logic_vector((3 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000",
    "000");
  signal op_mem_20_24_front_din: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((3 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0ca3374762 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0ca3374762;


architecture behavior of delay_0ca3374762 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (512 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(511);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 511 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_f1ac4bddff is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_f1ac4bddff;


architecture behavior of constant_f1ac4bddff is
begin
  op <= "0000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_498bc68c14 is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_498bc68c14;


architecture behavior of constant_498bc68c14 is
begin
  op <= "0000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fbc2f0cce1 is
  port (
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fbc2f0cce1;


architecture behavior of constant_fbc2f0cce1 is
begin
  op <= "1000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_d3720c25c3 is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((10 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_d3720c25c3;


architecture behavior of counter_d3720c25c3 is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((10 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((10 - 1) downto 0);
  signal count_reg_20_23: unsigned((10 - 1) downto 0) := "0000000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((12 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((12 - 1) downto 0);
  signal count_reg_join_48_3: signed((12 - 1) downto 0);
  signal count_reg_join_44_1: signed((12 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((10 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 12, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("000000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 12, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 10, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_0ffd72e037 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_0ffd72e037;


architecture behavior of relational_0ffd72e037 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_f6702ea2f7 is
  port (
    a : in std_logic_vector((10 - 1) downto 0);
    b : in std_logic_vector((10 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_f6702ea2f7;


architecture behavior of relational_f6702ea2f7 is
  signal a_1_31: unsigned((10 - 1) downto 0);
  signal b_1_34: unsigned((10 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_61242a554d is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_61242a554d;


architecture behavior of counter_61242a554d is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((10 - 1) downto 0) := "0000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((11 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("0000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_cf540617d5 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_cf540617d5;


architecture behavior of concat_cf540617d5 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_8f12c32de0 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_8f12c32de0;


architecture behavior of concat_8f12c32de0 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4ca77626c8 is
  port (
    d : in std_logic_vector((4 - 1) downto 0);
    q : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4ca77626c8;


architecture behavior of delay_4ca77626c8 is
  signal d_1_22: std_logic_vector((4 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000");
  signal op_mem_20_24_front_din: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_4f82bd00e5 is
  port (
    d : in std_logic_vector((4 - 1) downto 0);
    q : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_4f82bd00e5;


architecture behavior of delay_4f82bd00e5 is
  signal d_1_22: std_logic_vector((4 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000",
    "0000");
  signal op_mem_20_24_front_din: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((4 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_1f855d073b is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_1f855d073b;


architecture behavior of delay_1f855d073b is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (256 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(255);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 255 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b4ec9de7d1 is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b4ec9de7d1;


architecture behavior of constant_b4ec9de7d1 is
begin
  op <= "000000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd85eb7067 is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd85eb7067;


architecture behavior of constant_fd85eb7067 is
begin
  op <= "000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4a391b9a0e is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4a391b9a0e;


architecture behavior of constant_4a391b9a0e is
begin
  op <= "100000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_1dea202a2f is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((9 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_1dea202a2f;


architecture behavior of counter_1dea202a2f is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((9 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((9 - 1) downto 0);
  signal count_reg_20_23: unsigned((9 - 1) downto 0) := "000000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((11 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((11 - 1) downto 0);
  signal count_reg_join_48_3: signed((11 - 1) downto 0);
  signal count_reg_join_44_1: signed((11 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((9 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 11, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("00000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 11, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 9, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6c3ee657fa is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6c3ee657fa;


architecture behavior of relational_6c3ee657fa is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_78eac2928d is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_78eac2928d;


architecture behavior of relational_78eac2928d is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_d5d467f1b8 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_d5d467f1b8;


architecture behavior of counter_d5d467f1b8 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((9 - 1) downto 0) := "000000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((10 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2b3acb49f4 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2b3acb49f4;


architecture behavior of concat_2b3acb49f4 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((5 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ac785d9b37 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ac785d9b37;


architecture behavior of concat_ac785d9b37 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_ae3f02567e is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_ae3f02567e;


architecture behavior of concat_ae3f02567e is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_b096bcf164 is
  port (
    d : in std_logic_vector((5 - 1) downto 0);
    q : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_b096bcf164;


architecture behavior of delay_b096bcf164 is
  signal d_1_22: std_logic_vector((5 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000");
  signal op_mem_20_24_front_din: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_38f665f8aa is
  port (
    d : in std_logic_vector((5 - 1) downto 0);
    q : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_38f665f8aa;


architecture behavior of delay_38f665f8aa is
  signal d_1_22: std_logic_vector((5 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "00000",
    "00000");
  signal op_mem_20_24_front_din: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((5 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_c33e9b879a is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_c33e9b879a;


architecture behavior of delay_c33e9b879a is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (128 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(127);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 127 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_b437b02512 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_b437b02512;


architecture behavior of constant_b437b02512 is
begin
  op <= "00000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_91ef1678ca is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_91ef1678ca;


architecture behavior of constant_91ef1678ca is
begin
  op <= "00000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8aae5d3bb is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8aae5d3bb;


architecture behavior of constant_e8aae5d3bb is
begin
  op <= "10000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_a98fb09579 is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((8 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_a98fb09579;


architecture behavior of counter_a98fb09579 is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((8 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((8 - 1) downto 0);
  signal count_reg_20_23: unsigned((8 - 1) downto 0) := "00000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((10 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((10 - 1) downto 0);
  signal count_reg_join_48_3: signed((10 - 1) downto 0);
  signal count_reg_join_44_1: signed((10 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((8 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 10, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("0000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 10, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 8, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_54048c8b02 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54048c8b02;


architecture behavior of relational_54048c8b02 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_16235eb2bf is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_16235eb2bf;


architecture behavior of relational_16235eb2bf is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_11ccef49a2 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_11ccef49a2;


architecture behavior of counter_11ccef49a2 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((8 - 1) downto 0) := "00000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((9 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "00000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("00000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_2dc093ca7a is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_2dc093ca7a;


architecture behavior of concat_2dc093ca7a is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((6 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c6a9b6687e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c6a9b6687e;


architecture behavior of concat_c6a9b6687e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_75261c7c53 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_75261c7c53;


architecture behavior of concat_75261c7c53 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((5 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0b18d34058 is
  port (
    d : in std_logic_vector((6 - 1) downto 0);
    q : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0b18d34058;


architecture behavior of delay_0b18d34058 is
  signal d_1_22: std_logic_vector((6 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "000000");
  signal op_mem_20_24_front_din: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_da3bb0b159 is
  port (
    d : in std_logic_vector((6 - 1) downto 0);
    q : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_da3bb0b159;


architecture behavior of delay_da3bb0b159 is
  signal d_1_22: std_logic_vector((6 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000",
    "000000");
  signal op_mem_20_24_front_din: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((6 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_9b6c7a899e is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_9b6c7a899e;


architecture behavior of delay_9b6c7a899e is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (64 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(63);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 63 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_180df391de is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_180df391de;


architecture behavior of constant_180df391de is
begin
  op <= "0000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7244cd602b is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7244cd602b;


architecture behavior of constant_7244cd602b is
begin
  op <= "0000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7b07120b87 is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7b07120b87;


architecture behavior of constant_7b07120b87 is
begin
  op <= "1000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_82d8714dde is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((7 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_82d8714dde;


architecture behavior of counter_82d8714dde is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((7 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((7 - 1) downto 0);
  signal count_reg_20_23: unsigned((7 - 1) downto 0) := "0000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((9 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((9 - 1) downto 0);
  signal count_reg_join_48_3: signed((9 - 1) downto 0);
  signal count_reg_join_44_1: signed((9 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((7 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 9, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("000000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 9, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 7, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9a3978c602 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9a3978c602;


architecture behavior of relational_9a3978c602 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_23065a6aa3 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_23065a6aa3;


architecture behavior of relational_23065a6aa3 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_aaa565147f is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_aaa565147f;


architecture behavior of counter_aaa565147f is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((7 - 1) downto 0) := "0000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((8 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("0000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_eb5f1ca7f9 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_eb5f1ca7f9;


architecture behavior of concat_eb5f1ca7f9 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_83e473517e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_83e473517e;


architecture behavior of concat_83e473517e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((7 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_dc245eb1d2 is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_dc245eb1d2;


architecture behavior of concat_dc245eb1d2 is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_9066adfc41 is
  port (
    d : in std_logic_vector((7 - 1) downto 0);
    q : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_9066adfc41;


architecture behavior of delay_9066adfc41 is
  signal d_1_22: std_logic_vector((7 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "0000000");
  signal op_mem_20_24_front_din: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_8a9e828e57 is
  port (
    d : in std_logic_vector((7 - 1) downto 0);
    q : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_8a9e828e57;


architecture behavior of delay_8a9e828e57 is
  signal d_1_22: std_logic_vector((7 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "0000000",
    "0000000");
  signal op_mem_20_24_front_din: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((7 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_895e998e80 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_895e998e80;


architecture behavior of delay_895e998e80 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (32 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(31);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 31 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a267c870be is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a267c870be;


architecture behavior of constant_a267c870be is
begin
  op <= "000001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7ea0f2fff7 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7ea0f2fff7;


architecture behavior of constant_7ea0f2fff7 is
begin
  op <= "000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_961b61f8a1 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_961b61f8a1;


architecture behavior of constant_961b61f8a1 is
begin
  op <= "100000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_9686286f74 is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((6 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_9686286f74;


architecture behavior of counter_9686286f74 is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((6 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((6 - 1) downto 0);
  signal count_reg_20_23: unsigned((6 - 1) downto 0) := "000000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((8 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((8 - 1) downto 0);
  signal count_reg_join_48_3: signed((8 - 1) downto 0);
  signal count_reg_join_44_1: signed((8 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((6 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 8, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("00000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 8, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 6, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_931d61fb72 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_931d61fb72;


architecture behavior of relational_931d61fb72 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_fe487ce1c7 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_fe487ce1c7;


architecture behavior of relational_fe487ce1c7 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_7888581f80 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_7888581f80;


architecture behavior of counter_7888581f80 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((6 - 1) downto 0) := "000000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((7 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "000000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("000001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7673b9b993 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7673b9b993;


architecture behavior of concat_7673b9b993 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_1ece14600f is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_1ece14600f;


architecture behavior of concat_1ece14600f is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_f62149b02a is
  port (
    in0 : in std_logic_vector((2 - 1) downto 0);
    in1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_f62149b02a;


architecture behavior of concat_f62149b02a is
  signal in0_1_23: unsigned((2 - 1) downto 0);
  signal in1_1_27: unsigned((7 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_ebec135d8a is
  port (
    d : in std_logic_vector((8 - 1) downto 0);
    q : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_ebec135d8a;


architecture behavior of delay_ebec135d8a is
  signal d_1_22: std_logic_vector((8 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (1 - 1)) of std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    0 => "00000000");
  signal op_mem_20_24_front_din: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(0);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_23f848c85b is
  port (
    d : in std_logic_vector((8 - 1) downto 0);
    q : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_23f848c85b;


architecture behavior of delay_23f848c85b is
  signal d_1_22: std_logic_vector((8 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (2 - 1)) of std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "00000000",
    "00000000");
  signal op_mem_20_24_front_din: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((8 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(1);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 1 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_3a3620b5a6 is
  port (
    d : in std_logic_vector((36 - 1) downto 0);
    q : out std_logic_vector((36 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_3a3620b5a6;


architecture behavior of delay_3a3620b5a6 is
  signal d_1_22: std_logic_vector((36 - 1) downto 0);
  type array_type_op_mem_20_24 is array (0 to (16 - 1)) of std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24: array_type_op_mem_20_24 := (
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000",
    "000000000000000000000000000000000000");
  signal op_mem_20_24_front_din: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_back: std_logic_vector((36 - 1) downto 0);
  signal op_mem_20_24_push_front_pop_back_en: std_logic;
begin
  d_1_22 <= d;
  op_mem_20_24_back <= op_mem_20_24(15);
  proc_op_mem_20_24: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_20_24_push_front_pop_back_en = '1')) then
        for i in 15 downto 1 loop 
          op_mem_20_24(i) <= op_mem_20_24(i-1);
        end loop;
        op_mem_20_24(0) <= op_mem_20_24_front_din;
      end if;
    end if;
  end process proc_op_mem_20_24;
  op_mem_20_24_front_din <= d_1_22;
  op_mem_20_24_push_front_pop_back_en <= '1';
  q <= op_mem_20_24_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_582a3706dd is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_582a3706dd;


architecture behavior of constant_582a3706dd is
begin
  op <= "00001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fe72737ca0 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fe72737ca0;


architecture behavior of constant_fe72737ca0 is
begin
  op <= "00000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_ef0e2e5fc6 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_ef0e2e5fc6;


architecture behavior of constant_ef0e2e5fc6 is
begin
  op <= "10000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_9e5adb68be is
  port (
    load : in std_logic_vector((1 - 1) downto 0);
    din : in std_logic_vector((5 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_9e5adb68be;


architecture behavior of counter_9e5adb68be is
  signal load_1_29: boolean;
  signal din_1_35: unsigned((5 - 1) downto 0);
  signal en_1_45: boolean;
  signal count_reg_20_23_next: unsigned((5 - 1) downto 0);
  signal count_reg_20_23: unsigned((5 - 1) downto 0) := "00000";
  signal count_reg_20_23_en: std_logic;
  signal cast_54_19: signed((7 - 1) downto 0);
  signal count_reg_54_7_addsub: signed((7 - 1) downto 0);
  signal count_reg_join_48_3: signed((7 - 1) downto 0);
  signal count_reg_join_44_1: signed((7 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal cast_count_reg_20_23_next: unsigned((5 - 1) downto 0);
begin
  load_1_29 <= ((load) = "1");
  din_1_35 <= std_logic_vector_to_unsigned(din);
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23_next;
      end if;
    end if;
  end process proc_count_reg_20_23;
  cast_54_19 <= u2s_cast(count_reg_20_23, 0, 7, 0);
  count_reg_54_7_addsub <= cast_54_19 - std_logic_vector_to_signed("0000001");
  proc_if_48_3: process (count_reg_54_7_addsub, din_1_35, load_1_29)
  is
  begin
    if load_1_29 then
      count_reg_join_48_3 <= u2s_cast(din_1_35, 0, 7, 0);
    else 
      count_reg_join_48_3 <= count_reg_54_7_addsub;
    end if;
  end process proc_if_48_3;
  proc_if_44_1: process (count_reg_join_48_3, en_1_45)
  is
  begin
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else 
      count_reg_join_44_1_en <= '0';
    end if;
    count_reg_join_44_1 <= count_reg_join_48_3;
  end process proc_if_44_1;
  cast_count_reg_20_23_next <= s2u_cast(count_reg_join_44_1, 0, 5, 0);
  count_reg_20_23_next <= cast_count_reg_20_23_next;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9ece3c8c4e is
  port (
    a : in std_logic_vector((5 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9ece3c8c4e;


architecture behavior of relational_9ece3c8c4e is
  signal a_1_31: unsigned((5 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_dc5bc996c9 is
  port (
    a : in std_logic_vector((5 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_dc5bc996c9;


architecture behavior of relational_dc5bc996c9 is
  signal a_1_31: unsigned((5 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_743b50abe9 is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_743b50abe9;


architecture behavior of counter_743b50abe9 is
  signal rst_1_40: boolean;
  signal count_reg_20_23: unsigned((5 - 1) downto 0) := "00000";
  signal count_reg_20_23_rst: std_logic;
  signal bool_44_4: boolean;
  signal count_reg_join_44_1: unsigned((6 - 1) downto 0);
  signal count_reg_join_44_1_rst: std_logic;
  signal rst_limit_join_44_1: boolean;
begin
  rst_1_40 <= ((rst) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "00000";
      elsif (ce = '1') then 
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("00001");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    else 
      count_reg_join_44_1_rst <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    else 
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/delay0"

entity delay0_entity_f75f886771 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_f75f886771;

architecture structural of delay0_entity_f75f886771 is
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant_op_net: std_logic;
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal ram_data_out_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  reinterpret_out_output_port_net_x0 <= din;
  dout <= ram_data_out_net_x0;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter: entity work.counter_e110f0a1fc
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      op => counter_op_net
    );

  ram: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 36,
      core_name0 => "bmg_72_77dc1780892a0930",
      latency => 2
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      data_in => reinterpret_out_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => constant_op_net,
      data_out => ram_data_out_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/add_even_real/a_debus"

entity a_debus_entity_7fbb8fef33 is
  port (
    bus_in: in std_logic_vector(17 downto 0); 
    msb_lsb_out1: out std_logic_vector(17 downto 0)
  );
end a_debus_entity_7fbb8fef33;

architecture structural of a_debus_entity_7fbb8fef33 is
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x0 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 18,
      y_width => 18
    )
    port map (
      x => reinterpret2_output_port_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/add_even_real/op_bussify"

entity op_bussify_entity_ce6a4655d9 is
  port (
    in1: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(18 downto 0)
  );
end op_bussify_entity_ce6a4655d9;

architecture structural of op_bussify_entity_ce6a4655d9 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/add_even_real"

entity add_even_real_entity_0c9b1bec21 is
  port (
    a: in std_logic_vector(17 downto 0); 
    b: in std_logic_vector(17 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(18 downto 0)
  );
end add_even_real_entity_0c9b1bec21;

architecture structural of add_even_real_entity_0c9b1bec21 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x2: std_logic;
  signal clk_1_sg_x2: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x2 <= a;
  reinterpret2_output_port_net_x3 <= b;
  ce_1_sg_x2 <= ce_1;
  clk_1_sg_x2 <= clk_1;
  dout <= reinterpret1_output_port_net_x3;

  a_debus_7fbb8fef33: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret2_output_port_net_x2,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_59920783799a8e86",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x2,
      clk => clk_1_sg_x2,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  b_debus_10839fd766: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret2_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  op_bussify_ce6a4655d9: entity work.op_bussify_entity_ce6a4655d9
    port map (
      in1 => addsub1_s_net_x0,
      bus_out => reinterpret1_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_convert/bussify"

entity bussify_entity_904656ce6f is
  port (
    in1: in std_logic_vector(17 downto 0); 
    in2: in std_logic_vector(17 downto 0); 
    in3: in std_logic_vector(17 downto 0); 
    in4: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(71 downto 0)
  );
end bussify_entity_904656ce6f;

architecture structural of bussify_entity_904656ce6f is
  signal adder_s_net_x3: std_logic_vector(17 downto 0);
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(17 downto 0);

begin
  adder_s_net_x3 <= in1;
  adder_s_net_x4 <= in2;
  adder_s_net_x5 <= in3;
  adder_s_net_x6 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_a246e373e7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x3,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x4,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x5,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => adder_s_net_x6,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_convert/conv1"

entity conv1_entity_b7bb9c0ff9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(18 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end conv1_entity_b7bb9c0ff9;

architecture structural of conv1_entity_b7bb9c0ff9 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x4: std_logic;
  signal clk_1_sg_x4: std_logic;
  signal concat_y_net: std_logic_vector(19 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(19 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(18 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x4 <= ce_1;
  clk_1_sg_x4 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 19,
      a_width => 20,
      b_arith => xlUnsigned,
      b_bin_pt => 19,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 21,
      core_name0 => "addsb_11_0_ff0037ba5117ccc6",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 21,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 18
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      en => "1",
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 19,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_504cae28bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_convert/debus"

entity debus_entity_9e67f505ae is
  port (
    bus_in: in std_logic_vector(75 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out4: out std_logic_vector(18 downto 0); 
    out2: out std_logic_vector(18 downto 0); 
    out3: out std_logic_vector(18 downto 0)
  );
end debus_entity_9e67f505ae;

architecture structural of debus_entity_9e67f505ae is
  signal concatenate_y_net_x0: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);
  signal slice3_y_net: std_logic_vector(18 downto 0);
  signal slice4_y_net: std_logic_vector(18 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x1;
  msb_out4 <= reinterpret4_output_port_net_x1;
  out2 <= reinterpret2_output_port_net_x1;
  out3 <= reinterpret3_output_port_net_x1;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x1
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x1
    );

  reinterpret3: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x1
    );

  reinterpret4: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 38,
      new_msb => 56,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 57,
      new_msb => 75,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_convert"

entity bus_convert_entity_2e4c080be1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(71 downto 0)
  );
end bus_convert_entity_2e4c080be1;

architecture structural of bus_convert_entity_2e4c080be1 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal ce_1_sg_x8: std_logic;
  signal clk_1_sg_x8: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x8 <= ce_1;
  clk_1_sg_x8 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_904656ce6f: entity work.bussify_entity_904656ce6f
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_b7bb9c0ff9: entity work.conv1_entity_b7bb9c0ff9
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_da7fbfe370: entity work.conv1_entity_b7bb9c0ff9
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_6816298181: entity work.conv1_entity_b7bb9c0ff9
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_a2a5c12894: entity work.conv1_entity_b7bb9c0ff9
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_9e67f505ae: entity work.debus_entity_9e67f505ae
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_expand"

entity bus_expand_entity_56e25b700f is
  port (
    bus_in: in std_logic_vector(71 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out4: out std_logic_vector(17 downto 0); 
    out2: out std_logic_vector(17 downto 0); 
    out3: out std_logic_vector(17 downto 0)
  );
end bus_expand_entity_56e25b700f;

architecture structural of bus_expand_entity_56e25b700f is
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);
  signal slice3_y_net: std_logic_vector(17 downto 0);
  signal slice4_y_net: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x4 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 53,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 54,
      new_msb => 71,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x4,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_expand_a"

entity bus_expand_a_entity_b94579d477 is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out2: out std_logic_vector(17 downto 0)
  );
end bus_expand_a_entity_b94579d477;

architecture structural of bus_expand_a_entity_b94579d477 is
  signal reinterpret1_output_port_net_x6: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);

begin
  reinterpret_out_output_port_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x6;
  msb_out2 <= reinterpret2_output_port_net_x3;

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x6
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x3
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret_out_output_port_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => reinterpret_out_output_port_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_scale/bussify"

entity bussify_entity_a4c627ef16 is
  port (
    in1: in std_logic_vector(18 downto 0); 
    in2: in std_logic_vector(18 downto 0); 
    in3: in std_logic_vector(18 downto 0); 
    in4: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(75 downto 0)
  );
end bussify_entity_a4c627ef16;

architecture structural of bussify_entity_a4c627ef16 is
  signal concatenate_y_net_x3: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(18 downto 0);
  signal scale1_op_net_x0: std_logic_vector(18 downto 0);
  signal scale2_op_net_x0: std_logic_vector(18 downto 0);
  signal scale3_op_net_x0: std_logic_vector(18 downto 0);
  signal scale4_op_net_x0: std_logic_vector(18 downto 0);

begin
  scale1_op_net_x0 <= in1;
  scale2_op_net_x0 <= in2;
  scale3_op_net_x0 <= in3;
  scale4_op_net_x0 <= in4;
  bus_out <= concatenate_y_net_x3;

  concatenate: entity work.concat_2aea51ccde
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x3
    );

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale1_op_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale2_op_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale3_op_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => scale4_op_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_scale/debus"

entity debus_entity_b713d0483e is
  port (
    bus_in: in std_logic_vector(75 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out4: out std_logic_vector(18 downto 0); 
    out2: out std_logic_vector(18 downto 0); 
    out3: out std_logic_vector(18 downto 0)
  );
end debus_entity_b713d0483e;

architecture structural of debus_entity_b713d0483e is
  signal concat_y_net_x0: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);
  signal slice3_y_net: std_logic_vector(18 downto 0);
  signal slice4_y_net: std_logic_vector(18 downto 0);

begin
  concat_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 38,
      new_msb => 56,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 57,
      new_msb => 75,
      x_width => 76,
      y_width => 19
    )
    port map (
      x => concat_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/bus_scale"

entity bus_scale_entity_316a2a993e is
  port (
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(75 downto 0)
  );
end bus_scale_entity_316a2a993e;

architecture structural of bus_scale_entity_316a2a993e is
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(75 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal scale1_op_net_x0: std_logic_vector(18 downto 0);
  signal scale2_op_net_x0: std_logic_vector(18 downto 0);
  signal scale3_op_net_x0: std_logic_vector(18 downto 0);
  signal scale4_op_net_x0: std_logic_vector(18 downto 0);

begin
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x4;

  bussify_a4c627ef16: entity work.bussify_entity_a4c627ef16
    port map (
      in1 => scale1_op_net_x0,
      in2 => scale2_op_net_x0,
      in3 => scale3_op_net_x0,
      in4 => scale4_op_net_x0,
      bus_out => concatenate_y_net_x4
    );

  debus_b713d0483e: entity work.debus_entity_b713d0483e
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  scale1: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret4_output_port_net_x0,
      op => scale1_op_net_x0
    );

  scale2: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret3_output_port_net_x0,
      op => scale2_op_net_x0
    );

  scale3: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret2_output_port_net_x0,
      op => scale3_op_net_x0
    );

  scale4: entity work.scale_9f61027ba4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret1_output_port_net_x0,
      op => scale4_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/munge_a/join"

entity join_entity_92d8cf050f is
  port (
    in1: in std_logic_vector(17 downto 0); 
    in2: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end join_entity_92d8cf050f;

architecture structural of join_entity_92d8cf050f is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x1 <= in1;
  reinterpret1_output_port_net_x1 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret1_output_port_net_x1,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/munge_a"

entity munge_a_entity_7fbc079bee is
  port (
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end munge_a_entity_7fbc079bee;

architecture structural of munge_a_entity_7fbc079bee is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal mux0_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(35 downto 0);

begin
  mux0_y_net_x0 <= din;
  dout <= reinterpret_out_output_port_net_x1;

  join_92d8cf050f: entity work.join_entity_92d8cf050f
    port map (
      in1 => reinterpret2_output_port_net_x2,
      in2 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x0
    );

  reinterpret: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux0_y_net_x0,
      output_port => reinterpret_output_port_net_x0
    );

  reinterpret_out: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x0,
      output_port => reinterpret_out_output_port_net_x1
    );

  split_04aa63b12a: entity work.bus_expand_a_entity_b94579d477
    port map (
      bus_in => reinterpret_output_port_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/ri_to_c"

entity ri_to_c_entity_5ed1c1a8f6 is
  port (
    im: in std_logic_vector(17 downto 0); 
    re: in std_logic_vector(17 downto 0); 
    c: out std_logic_vector(35 downto 0)
  );
end ri_to_c_entity_5ed1c1a8f6;

architecture structural of ri_to_c_entity_5ed1c1a8f6 is
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal force_im_output_port_net: std_logic_vector(17 downto 0);
  signal force_re_output_port_net: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  reinterpret2_output_port_net_x1 <= im;
  reinterpret4_output_port_net_x1 <= re;
  c <= concat_y_net_x1;

  concat: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x1
    );

  force_im: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_9306b5127f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x1,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0/sub_even_imag"

entity sub_even_imag_entity_27636760b6 is
  port (
    a: in std_logic_vector(17 downto 0); 
    b: in std_logic_vector(17 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(18 downto 0)
  );
end sub_even_imag_entity_27636760b6;

architecture structural of sub_even_imag_entity_27636760b6 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x9: std_logic;
  signal clk_1_sg_x9: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x12: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(17 downto 0);

begin
  reinterpret1_output_port_net_x11 <= a;
  reinterpret1_output_port_net_x12 <= b;
  ce_1_sg_x9 <= ce_1;
  clk_1_sg_x9 <= clk_1;
  dout <= reinterpret1_output_port_net_x13;

  a_debus_9c22b08e03: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret1_output_port_net_x11,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_18f6f1cec46d694e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x9,
      ce => ce_1_sg_x9,
      clk => clk_1_sg_x9,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  b_debus_8079305c23: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret1_output_port_net_x12,
      msb_lsb_out1 => reinterpret1_output_port_net_x9
    );

  op_bussify_835cfde070: entity work.op_bussify_entity_ce6a4655d9
    port map (
      in1 => addsub1_s_net_x0,
      bus_out => reinterpret1_output_port_net_x13
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/hilbert0"

entity hilbert0_entity_99acf82149 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    even: out std_logic_vector(35 downto 0); 
    odd: out std_logic_vector(35 downto 0)
  );
end hilbert0_entity_99acf82149;

architecture structural of hilbert0_entity_99acf82149 is
  signal ce_1_sg_x11: std_logic;
  signal clk_1_sg_x11: std_logic;
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concat_y_net_x2: std_logic_vector(35 downto 0);
  signal concat_y_net_x3: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(75 downto 0);
  signal mux0_y_net_x1: std_logic_vector(35 downto 0);
  signal mux1_y_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x12: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);

begin
  mux0_y_net_x1 <= a;
  mux1_y_net_x1 <= b;
  ce_1_sg_x11 <= ce_1;
  clk_1_sg_x11 <= clk_1;
  even <= reinterpret_out_output_port_net_x5;
  odd <= reinterpret_out_output_port_net_x6;

  add_even_real_0c9b1bec21: entity work.add_even_real_entity_0c9b1bec21
    port map (
      a => reinterpret2_output_port_net_x6,
      b => reinterpret2_output_port_net_x7,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x3
    );

  add_odd_real_1857588202: entity work.add_even_real_entity_0c9b1bec21
    port map (
      a => reinterpret1_output_port_net_x11,
      b => reinterpret1_output_port_net_x12,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x7
    );

  bus_convert_2e4c080be1: entity work.bus_convert_entity_2e4c080be1
    port map (
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      din => concatenate_y_net_x5,
      dout => concatenate_y_net_x4
    );

  bus_expand_56e25b700f: entity work.bus_expand_entity_56e25b700f
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

  bus_expand_a_b94579d477: entity work.bus_expand_a_entity_b94579d477
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => reinterpret2_output_port_net_x6
    );

  bus_expand_b_258073bd02: entity work.bus_expand_a_entity_b94579d477
    port map (
      bus_in => reinterpret_out_output_port_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x12,
      msb_out2 => reinterpret2_output_port_net_x7
    );

  bus_scale_316a2a993e: entity work.bus_scale_entity_316a2a993e
    port map (
      din => concat_y_net_x1,
      dout => concatenate_y_net_x5
    );

  concat: entity work.concat_2aea51ccde
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net_x3,
      in1 => reinterpret1_output_port_net_x4,
      in2 => reinterpret1_output_port_net_x13,
      in3 => reinterpret1_output_port_net_x7,
      y => concat_y_net_x1
    );

  munge_a_7fbc079bee: entity work.munge_a_entity_7fbc079bee
    port map (
      din => mux0_y_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_b_fc82ab8c7f: entity work.munge_a_entity_7fbc079bee
    port map (
      din => mux1_y_net_x1,
      dout => reinterpret_out_output_port_net_x2
    );

  munge_even_f72c5aa202: entity work.munge_a_entity_7fbc079bee
    port map (
      din => concat_y_net_x2,
      dout => reinterpret_out_output_port_net_x5
    );

  munge_odd_5045b10a0c: entity work.munge_a_entity_7fbc079bee
    port map (
      din => concat_y_net_x3,
      dout => reinterpret_out_output_port_net_x6
    );

  ri_to_c1_353b44a8e3: entity work.ri_to_c_entity_5ed1c1a8f6
    port map (
      im => reinterpret3_output_port_net_x1,
      re => reinterpret1_output_port_net_x1,
      c => concat_y_net_x3
    );

  ri_to_c_5ed1c1a8f6: entity work.ri_to_c_entity_5ed1c1a8f6
    port map (
      im => reinterpret2_output_port_net_x1,
      re => reinterpret4_output_port_net_x1,
      c => concat_y_net_x2
    );

  sub_even_imag_27636760b6: entity work.sub_even_imag_entity_27636760b6
    port map (
      a => reinterpret1_output_port_net_x11,
      b => reinterpret1_output_port_net_x12,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x13
    );

  sub_odd_imag_9979230f77: entity work.sub_even_imag_entity_27636760b6
    port map (
      a => reinterpret2_output_port_net_x7,
      b => reinterpret2_output_port_net_x6,
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      dout => reinterpret1_output_port_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/complex_conj0/imag_negate/bussify"

entity bussify_entity_7962d3f7d8 is
  port (
    in1: in std_logic_vector(17 downto 0); 
    bus_out: out std_logic_vector(17 downto 0)
  );
end bussify_entity_7962d3f7d8;

architecture structural of bussify_entity_7962d3f7d8 is
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);

begin
  neg1_op_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => neg1_op_net_x0,
      output_port => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/complex_conj0/imag_negate"

entity imag_negate_entity_89e12f4fc9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(17 downto 0); 
    dout: out std_logic_vector(17 downto 0)
  );
end imag_negate_entity_89e12f4fc9;

architecture structural of imag_negate_entity_89e12f4fc9 is
  signal ce_1_sg_x22: std_logic;
  signal clk_1_sg_x22: std_logic;
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x22 <= ce_1;
  clk_1_sg_x22 <= clk_1;
  reinterpret1_output_port_net_x4 <= din;
  dout <= reinterpret1_output_port_net_x5;

  bussify_7962d3f7d8: entity work.bussify_entity_7962d3f7d8
    port map (
      in1 => neg1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x5
    );

  debus_5788bba85e: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret1_output_port_net_x4,
      msb_lsb_out1 => reinterpret1_output_port_net_x3
    );

  neg1: entity work.negate_f983e30a8b
    port map (
      ce => ce_1_sg_x22,
      clk => clk_1_sg_x22,
      clr => '0',
      ip => reinterpret1_output_port_net_x3,
      op => neg1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/complex_conj0"

entity complex_conj0_entity_e5a1b463f3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    z: in std_logic_vector(35 downto 0); 
    z_x0: out std_logic_vector(35 downto 0)
  );
end complex_conj0_entity_e5a1b463f3;

architecture structural of complex_conj0_entity_e5a1b463f3 is
  signal ce_1_sg_x23: std_logic;
  signal clk_1_sg_x23: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal d3_q_net_x1: std_logic_vector(35 downto 0);
  signal real_delay_q_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x23 <= ce_1;
  clk_1_sg_x23 <= clk_1;
  d3_q_net_x1 <= z;
  z_x0 <= reinterpret_out_output_port_net_x2;

  bus_create_f1bd892860: entity work.join_entity_92d8cf050f
    port map (
      in1 => real_delay_q_net_x0,
      in2 => reinterpret1_output_port_net_x5,
      bus_out => concatenate_y_net_x2
    );

  bus_expand_41a2a65fe0: entity work.bus_expand_a_entity_b94579d477
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  imag_negate_89e12f4fc9: entity work.imag_negate_entity_89e12f4fc9
    port map (
      ce_1 => ce_1_sg_x23,
      clk_1 => clk_1_sg_x23,
      din => reinterpret1_output_port_net_x4,
      dout => reinterpret1_output_port_net_x5
    );

  munge_in_a6fb6151c7: entity work.munge_a_entity_7fbc079bee
    port map (
      din => d3_q_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_out_24928d72f4: entity work.munge_a_entity_7fbc079bee
    port map (
      din => concatenate_y_net_x2,
      dout => reinterpret_out_output_port_net_x2
    );

  real_delay: entity work.delay_6699ee0916
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x0,
      q => real_delay_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/dmux0/d_bussify"

entity d_bussify_entity_edab46ac75 is
  port (
    in1: in std_logic_vector(35 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end d_bussify_entity_edab46ac75;

architecture structural of d_bussify_entity_edab46ac75 is
  signal mux0_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);

begin
  mux0_y_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux0_y_net_x0,
      output_port => reinterpret1_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/dmux0/expand0"

entity expand0_entity_49f6172f66 is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    msb_lsb_out1: out std_logic_vector(35 downto 0)
  );
end expand0_entity_49f6172f66;

architecture structural of expand0_entity_49f6172f66 is
  signal delay0_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);

begin
  delay0_q_net_x0 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 36,
      y_width => 36
    )
    port map (
      x => delay0_q_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/dmux0/sel_expand"

entity sel_expand_entity_894fe05a71 is
  port (
    bus_in: in std_logic; 
    msb_lsb_out1: out std_logic
  );
end sel_expand_entity_894fe05a71;

architecture structural of sel_expand_entity_894fe05a71 is
  signal reinterpret1_output_port_net_x1: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic;
  signal slice1_y_net: std_logic;

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_81130c7f2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => slice1_y_net,
      output_port(0) => reinterpret1_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 1,
      y_width => 1
    )
    port map (
      x(0) => reinterpret1_output_port_net_x1,
      y(0) => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/dmux0"

entity dmux0_entity_5714570cb6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d0: in std_logic_vector(35 downto 0); 
    d1: in std_logic_vector(35 downto 0); 
    sel: in std_logic; 
    out_x0: out std_logic_vector(35 downto 0)
  );
end dmux0_entity_5714570cb6;

architecture structural of dmux0_entity_5714570cb6 is
  signal ce_1_sg_x30: std_logic;
  signal clk_1_sg_x30: std_logic;
  signal delay0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux0_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic;
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x4: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x30 <= ce_1;
  clk_1_sg_x30 <= clk_1;
  delay0_q_net_x1 <= d0;
  reinterpret_out_output_port_net_x4 <= d1;
  reinterpret1_output_port_net_x5 <= sel;
  out_x0 <= reinterpret1_output_port_net_x6;

  d_bussify_edab46ac75: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => mux0_y_net_x0,
      bus_out => reinterpret1_output_port_net_x6
    );

  expand0_49f6172f66: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => delay0_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  expand1_1d738941cf: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret_out_output_port_net_x4,
      msb_lsb_out1 => reinterpret1_output_port_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      d0 => reinterpret1_output_port_net_x1,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => reinterpret1_output_port_net_x3,
      y => mux0_y_net_x0
    );

  sel_expand_894fe05a71: entity work.sel_expand_entity_894fe05a71
    port map (
      bus_in => reinterpret1_output_port_net_x5,
      msb_lsb_out1 => reinterpret1_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/sel_replicate0/bussify"

entity bussify_entity_ad099992fc is
  port (
    in1: in std_logic; 
    bus_out: out std_logic
  );
end bussify_entity_ad099992fc;

architecture structural of bussify_entity_ad099992fc is
  signal reinterpret1_output_port_net_x6: std_logic;
  signal relational_op_net_x0: std_logic;

begin
  relational_op_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x6;

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => relational_op_net_x0,
      output_port(0) => reinterpret1_output_port_net_x6
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum/sel_replicate0"

entity sel_replicate0_entity_bc92d7dfef is
  port (
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sel_replicate0_entity_bc92d7dfef;

architecture structural of sel_replicate0_entity_bc92d7dfef is
  signal reinterpret1_output_port_net_x7: std_logic;
  signal relational_op_net_x1: std_logic;

begin
  relational_op_net_x1 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x7;

  bussify_ad099992fc: entity work.bussify_entity_ad099992fc
    port map (
      in1 => relational_op_net_x1,
      bus_out => reinterpret1_output_port_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/mirror_spectrum"

entity mirror_spectrum_entity_dc7f261b12 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    din1: in std_logic_vector(35 downto 0); 
    din2: in std_logic_vector(35 downto 0); 
    din3: in std_logic_vector(35 downto 0); 
    reo_in0: in std_logic_vector(35 downto 0); 
    reo_in1: in std_logic_vector(35 downto 0); 
    reo_in2: in std_logic_vector(35 downto 0); 
    reo_in3: in std_logic_vector(35 downto 0); 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    dout1: out std_logic_vector(35 downto 0); 
    dout2: out std_logic_vector(35 downto 0); 
    dout3: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end mirror_spectrum_entity_dc7f261b12;

architecture structural of mirror_spectrum_entity_dc7f261b12 is
  signal ce_1_sg_x34: std_logic;
  signal clk_1_sg_x34: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal d3_q_net_x2: std_logic_vector(35 downto 0);
  signal d4_q_net_x2: std_logic_vector(35 downto 0);
  signal d5_q_net_x2: std_logic_vector(35 downto 0);
  signal d6_q_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net_x1: std_logic_vector(35 downto 0);
  signal delay1_q_net_x1: std_logic_vector(35 downto 0);
  signal delay2_q_net_x1: std_logic_vector(35 downto 0);
  signal delay3_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x0: std_logic;
  signal ram_data_out_net_x2: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic;
  signal reinterpret1_output_port_net_x12: std_logic;
  signal reinterpret1_output_port_net_x13: std_logic;
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x9: std_logic_vector(35 downto 0);
  signal relational_op_net_x7: std_logic;
  signal sync_delay0_q_net: std_logic;
  signal sync_delay1_q_net_x0: std_logic;

begin
  ce_1_sg_x34 <= ce_1;
  clk_1_sg_x34 <= clk_1;
  ram_data_out_net_x2 <= din0;
  ram_data_out_net_x3 <= din1;
  reinterpret_out_output_port_net_x10 <= din2;
  reinterpret_out_output_port_net_x11 <= din3;
  d3_q_net_x2 <= reo_in0;
  d4_q_net_x2 <= reo_in1;
  d5_q_net_x2 <= reo_in2;
  d6_q_net_x2 <= reo_in3;
  mux_y_net_x0 <= sync;
  dout0 <= reinterpret1_output_port_net_x14;
  dout1 <= reinterpret1_output_port_net_x15;
  dout2 <= reinterpret1_output_port_net_x16;
  dout3 <= reinterpret1_output_port_net_x17;
  sync_out <= sync_delay1_q_net_x0;

  complex_conj0_e5a1b463f3: entity work.complex_conj0_entity_e5a1b463f3
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      z => d3_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x6
    );

  complex_conj1_73a353caef: entity work.complex_conj0_entity_e5a1b463f3
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      z => d4_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x7
    );

  complex_conj2_5e819d55af: entity work.complex_conj0_entity_e5a1b463f3
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      z => d5_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x8
    );

  complex_conj3_a0ce88ea3d: entity work.complex_conj0_entity_e5a1b463f3
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      z => d6_q_net_x2,
      z_x0 => reinterpret_out_output_port_net_x9
    );

  constant_x0: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_c48d6dcab5
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      rst(0) => sync_delay0_q_net,
      op => counter_op_net
    );

  delay0: entity work.delay_6096a10519
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => ram_data_out_net_x2,
      q => delay0_q_net_x1
    );

  delay1: entity work.delay_6096a10519
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => ram_data_out_net_x3,
      q => delay1_q_net_x1
    );

  delay2: entity work.delay_6096a10519
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => reinterpret_out_output_port_net_x10,
      q => delay2_q_net_x1
    );

  delay3: entity work.delay_6096a10519
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d => reinterpret_out_output_port_net_x11,
      q => delay3_q_net_x1
    );

  dmux0_5714570cb6: entity work.dmux0_entity_5714570cb6
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      d0 => delay0_q_net_x1,
      d1 => reinterpret_out_output_port_net_x6,
      sel => reinterpret1_output_port_net_x10,
      out_x0 => reinterpret1_output_port_net_x14
    );

  dmux1_87e5c37770: entity work.dmux0_entity_5714570cb6
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      d0 => delay1_q_net_x1,
      d1 => reinterpret_out_output_port_net_x7,
      sel => reinterpret1_output_port_net_x11,
      out_x0 => reinterpret1_output_port_net_x15
    );

  dmux2_2b2adfca5d: entity work.dmux0_entity_5714570cb6
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      d0 => delay2_q_net_x1,
      d1 => reinterpret_out_output_port_net_x8,
      sel => reinterpret1_output_port_net_x12,
      out_x0 => reinterpret1_output_port_net_x16
    );

  dmux3_db6b9a62c4: entity work.dmux0_entity_5714570cb6
    port map (
      ce_1 => ce_1_sg_x34,
      clk_1 => clk_1_sg_x34,
      d0 => delay3_q_net_x1,
      d1 => reinterpret_out_output_port_net_x9,
      sel => reinterpret1_output_port_net_x13,
      out_x0 => reinterpret1_output_port_net_x17
    );

  relational: entity work.relational_54e7975215
    port map (
      a => counter_op_net,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net_x7
    );

  sel_replicate0_bc92d7dfef: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => relational_op_net_x7,
      out_x0 => reinterpret1_output_port_net_x10
    );

  sel_replicate1_9bc4511ef8: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => relational_op_net_x7,
      out_x0 => reinterpret1_output_port_net_x11
    );

  sel_replicate2_4c49384471: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => relational_op_net_x7,
      out_x0 => reinterpret1_output_port_net_x12
    );

  sel_replicate3_820f5d70e5: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => relational_op_net_x7,
      out_x0 => reinterpret1_output_port_net_x13
    );

  sync_delay0: entity work.delay_e055964d40
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => sync_delay0_q_net
    );

  sync_delay1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x34,
      clk => clk_1_sg_x34,
      clr => '0',
      d(0) => sync_delay0_q_net,
      q(0) => sync_delay1_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/addr_expand"

entity addr_expand_entity_8d8c5a295c is
  port (
    bus_in: in std_logic_vector(11 downto 0); 
    msb_lsb_out1: out std_logic_vector(11 downto 0)
  );
end addr_expand_entity_8d8c5a295c;

architecture structural of addr_expand_entity_8d8c5a295c is
  signal reinterpret1_output_port_net_x1: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(11 downto 0);
  signal slice1_y_net: std_logic_vector(11 downto 0);

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 12,
      y_width => 12
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/addr_replicate/bussify"

entity bussify_entity_9313117430 is
  port (
    in1: in std_logic_vector(11 downto 0); 
    bus_out: out std_logic_vector(11 downto 0)
  );
end bussify_entity_9313117430;

architecture structural of bussify_entity_9313117430 is
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(11 downto 0);

begin
  mux_y_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x0,
      output_port => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/addr_replicate"

entity addr_replicate_entity_cc9047aff8 is
  port (
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(11 downto 0)
  );
end addr_replicate_entity_cc9047aff8;

architecture structural of addr_replicate_entity_cc9047aff8 is
  signal mux_y_net_x1: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(11 downto 0);

begin
  mux_y_net_x1 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x3;

  bussify_9313117430: entity work.bussify_entity_9313117430
    port map (
      in1 => mux_y_net_x1,
      bus_out => reinterpret1_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/debus_addr"

entity debus_addr_entity_683e5a971d is
  port (
    bus_in: in std_logic_vector(107 downto 0); 
    lsb_out1: out std_logic_vector(11 downto 0); 
    msb_out9: out std_logic_vector(11 downto 0); 
    out2: out std_logic_vector(11 downto 0); 
    out3: out std_logic_vector(11 downto 0); 
    out4: out std_logic_vector(11 downto 0); 
    out5: out std_logic_vector(11 downto 0); 
    out6: out std_logic_vector(11 downto 0); 
    out7: out std_logic_vector(11 downto 0); 
    out8: out std_logic_vector(11 downto 0)
  );
end debus_addr_entity_683e5a971d;

architecture structural of debus_addr_entity_683e5a971d is
  signal concatenate_y_net_x0: std_logic_vector(107 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret5_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret6_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret7_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret8_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret9_output_port_net_x0: std_logic_vector(11 downto 0);
  signal slice1_y_net: std_logic_vector(11 downto 0);
  signal slice2_y_net: std_logic_vector(11 downto 0);
  signal slice3_y_net: std_logic_vector(11 downto 0);
  signal slice4_y_net: std_logic_vector(11 downto 0);
  signal slice5_y_net: std_logic_vector(11 downto 0);
  signal slice6_y_net: std_logic_vector(11 downto 0);
  signal slice7_y_net: std_logic_vector(11 downto 0);
  signal slice8_y_net: std_logic_vector(11 downto 0);
  signal slice9_y_net: std_logic_vector(11 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out9 <= reinterpret9_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;
  out4 <= reinterpret4_output_port_net_x0;
  out5 <= reinterpret5_output_port_net_x0;
  out6 <= reinterpret6_output_port_net_x0;
  out7 <= reinterpret7_output_port_net_x0;
  out8 <= reinterpret8_output_port_net_x0;

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  reinterpret5: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice5_y_net,
      output_port => reinterpret5_output_port_net_x0
    );

  reinterpret6: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice6_y_net,
      output_port => reinterpret6_output_port_net_x0
    );

  reinterpret7: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice7_y_net,
      output_port => reinterpret7_output_port_net_x0
    );

  reinterpret8: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice8_y_net,
      output_port => reinterpret8_output_port_net_x0
    );

  reinterpret9: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice9_y_net,
      output_port => reinterpret9_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 23,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 35,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 47,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

  slice5: entity work.xlslice
    generic map (
      new_lsb => 48,
      new_msb => 59,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice5_y_net
    );

  slice6: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 71,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice6_y_net
    );

  slice7: entity work.xlslice
    generic map (
      new_lsb => 72,
      new_msb => 83,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice7_y_net
    );

  slice8: entity work.xlslice
    generic map (
      new_lsb => 84,
      new_msb => 95,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice8_y_net
    );

  slice9: entity work.xlslice
    generic map (
      new_lsb => 96,
      new_msb => 107,
      x_width => 108,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice9_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/debus_din"

entity debus_din_entity_d2fe8dc95c is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(3 downto 0); 
    msb_out9: out std_logic_vector(3 downto 0); 
    out2: out std_logic_vector(3 downto 0); 
    out3: out std_logic_vector(3 downto 0); 
    out4: out std_logic_vector(3 downto 0); 
    out5: out std_logic_vector(3 downto 0); 
    out6: out std_logic_vector(3 downto 0); 
    out7: out std_logic_vector(3 downto 0); 
    out8: out std_logic_vector(3 downto 0)
  );
end debus_din_entity_d2fe8dc95c;

architecture structural of debus_din_entity_d2fe8dc95c is
  signal ddin_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret5_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret6_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret7_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret8_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret9_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net: std_logic_vector(3 downto 0);
  signal slice2_y_net: std_logic_vector(3 downto 0);
  signal slice3_y_net: std_logic_vector(3 downto 0);
  signal slice4_y_net: std_logic_vector(3 downto 0);
  signal slice5_y_net: std_logic_vector(3 downto 0);
  signal slice6_y_net: std_logic_vector(3 downto 0);
  signal slice7_y_net: std_logic_vector(3 downto 0);
  signal slice8_y_net: std_logic_vector(3 downto 0);
  signal slice9_y_net: std_logic_vector(3 downto 0);

begin
  ddin_q_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out9 <= reinterpret9_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;
  out4 <= reinterpret4_output_port_net_x0;
  out5 <= reinterpret5_output_port_net_x0;
  out6 <= reinterpret6_output_port_net_x0;
  out7 <= reinterpret7_output_port_net_x0;
  out8 <= reinterpret8_output_port_net_x0;

  reinterpret1: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  reinterpret5: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice5_y_net,
      output_port => reinterpret5_output_port_net_x0
    );

  reinterpret6: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice6_y_net,
      output_port => reinterpret6_output_port_net_x0
    );

  reinterpret7: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice7_y_net,
      output_port => reinterpret7_output_port_net_x0
    );

  reinterpret8: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice8_y_net,
      output_port => reinterpret8_output_port_net_x0
    );

  reinterpret9: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice9_y_net,
      output_port => reinterpret9_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 7,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 11,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 15,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice4_y_net
    );

  slice5: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 19,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice5_y_net
    );

  slice6: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 23,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice6_y_net
    );

  slice7: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 27,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice7_y_net
    );

  slice8: entity work.xlslice
    generic map (
      new_lsb => 28,
      new_msb => 31,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice8_y_net
    );

  slice9: entity work.xlslice
    generic map (
      new_lsb => 32,
      new_msb => 35,
      x_width => 36,
      y_width => 4
    )
    port map (
      x => ddin_q_net_x0,
      y => slice9_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/debus_we"

entity debus_we_entity_118daa2628 is
  port (
    bus_in: in std_logic_vector(8 downto 0); 
    lsb_out1: out std_logic; 
    msb_out9: out std_logic; 
    out2: out std_logic; 
    out3: out std_logic; 
    out4: out std_logic; 
    out5: out std_logic; 
    out6: out std_logic; 
    out7: out std_logic; 
    out8: out std_logic
  );
end debus_we_entity_118daa2628;

architecture structural of debus_we_entity_118daa2628 is
  signal concatenate_y_net_x0: std_logic_vector(8 downto 0);
  signal slice1_y_net_x0: std_logic;
  signal slice2_y_net_x0: std_logic;
  signal slice3_y_net_x0: std_logic;
  signal slice4_y_net_x0: std_logic;
  signal slice5_y_net_x0: std_logic;
  signal slice6_y_net_x0: std_logic;
  signal slice7_y_net_x0: std_logic;
  signal slice8_y_net_x0: std_logic;
  signal slice9_y_net_x0: std_logic;

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= slice1_y_net_x0;
  msb_out9 <= slice9_y_net_x0;
  out2 <= slice2_y_net_x0;
  out3 <= slice3_y_net_x0;
  out4 <= slice4_y_net_x0;
  out5 <= slice5_y_net_x0;
  out6 <= slice6_y_net_x0;
  out7 <= slice7_y_net_x0;
  out8 <= slice8_y_net_x0;

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice1_y_net_x0
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice2_y_net_x0
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice3_y_net_x0
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice4_y_net_x0
    );

  slice5: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice5_y_net_x0
    );

  slice6: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice6_y_net_x0
    );

  slice7: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice7_y_net_x0
    );

  slice8: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice8_y_net_x0
    );

  slice9: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice9_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/din_bussify"

entity din_bussify_entity_e936a8b4d0 is
  port (
    in1: in std_logic_vector(3 downto 0); 
    in2: in std_logic_vector(3 downto 0); 
    in3: in std_logic_vector(3 downto 0); 
    in4: in std_logic_vector(3 downto 0); 
    in5: in std_logic_vector(3 downto 0); 
    in6: in std_logic_vector(3 downto 0); 
    in7: in std_logic_vector(3 downto 0); 
    in8: in std_logic_vector(3 downto 0); 
    in9: in std_logic_vector(3 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end din_bussify_entity_e936a8b4d0;

architecture structural of din_bussify_entity_e936a8b4d0 is
  signal bram0_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram4_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram5_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram6_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram7_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram8_data_out_net_x0: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret5_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret6_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret7_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret8_output_port_net: std_logic_vector(3 downto 0);
  signal reinterpret9_output_port_net: std_logic_vector(3 downto 0);

begin
  bram0_data_out_net_x0 <= in1;
  bram1_data_out_net_x0 <= in2;
  bram2_data_out_net_x0 <= in3;
  bram3_data_out_net_x0 <= in4;
  bram4_data_out_net_x0 <= in5;
  bram5_data_out_net_x0 <= in6;
  bram6_data_out_net_x0 <= in7;
  bram7_data_out_net_x0 <= in8;
  bram8_data_out_net_x0 <= in9;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_e4837c85a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      in4 => reinterpret5_output_port_net,
      in5 => reinterpret6_output_port_net,
      in6 => reinterpret7_output_port_net,
      in7 => reinterpret8_output_port_net,
      in8 => reinterpret9_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram0_data_out_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram1_data_out_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram2_data_out_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram3_data_out_net_x0,
      output_port => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram4_data_out_net_x0,
      output_port => reinterpret5_output_port_net
    );

  reinterpret6: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram5_data_out_net_x0,
      output_port => reinterpret6_output_port_net
    );

  reinterpret7: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram6_data_out_net_x0,
      output_port => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram7_data_out_net_x0,
      output_port => reinterpret8_output_port_net
    );

  reinterpret9: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram8_data_out_net_x0,
      output_port => reinterpret9_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/rep_addr/bussify"

entity bussify_entity_8403f05c85 is
  port (
    in1: in std_logic_vector(11 downto 0); 
    in2: in std_logic_vector(11 downto 0); 
    in3: in std_logic_vector(11 downto 0); 
    in4: in std_logic_vector(11 downto 0); 
    in5: in std_logic_vector(11 downto 0); 
    in6: in std_logic_vector(11 downto 0); 
    in7: in std_logic_vector(11 downto 0); 
    in8: in std_logic_vector(11 downto 0); 
    in9: in std_logic_vector(11 downto 0); 
    bus_out: out std_logic_vector(107 downto 0)
  );
end bussify_entity_8403f05c85;

architecture structural of bussify_entity_8403f05c85 is
  signal concatenate_y_net_x1: std_logic_vector(107 downto 0);
  signal din3_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_2_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_3_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_4_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_5_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_6_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_7_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_8_q_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret5_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret6_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret7_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret8_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret9_output_port_net: std_logic_vector(11 downto 0);

begin
  din3_0_q_net_x0 <= in1;
  din3_1_q_net_x0 <= in2;
  din3_2_q_net_x0 <= in3;
  din3_3_q_net_x0 <= in4;
  din3_4_q_net_x0 <= in5;
  din3_5_q_net_x0 <= in6;
  din3_6_q_net_x0 <= in7;
  din3_7_q_net_x0 <= in8;
  din3_8_q_net_x0 <= in9;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_336ab7141a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      in4 => reinterpret5_output_port_net,
      in5 => reinterpret6_output_port_net,
      in6 => reinterpret7_output_port_net,
      in7 => reinterpret8_output_port_net,
      in8 => reinterpret9_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_0_q_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_1_q_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_2_q_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_3_q_net_x0,
      output_port => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_4_q_net_x0,
      output_port => reinterpret5_output_port_net
    );

  reinterpret6: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_5_q_net_x0,
      output_port => reinterpret6_output_port_net
    );

  reinterpret7: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_6_q_net_x0,
      output_port => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_7_q_net_x0,
      output_port => reinterpret8_output_port_net
    );

  reinterpret9: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_8_q_net_x0,
      output_port => reinterpret9_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/rep_addr"

entity rep_addr_entity_152c8d6b28 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(107 downto 0)
  );
end rep_addr_entity_152c8d6b28;

architecture structural of rep_addr_entity_152c8d6b28 is
  signal ce_1_sg_x35: std_logic;
  signal clk_1_sg_x35: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(107 downto 0);
  signal din0_0_q_net: std_logic_vector(11 downto 0);
  signal din1_0_q_net: std_logic_vector(11 downto 0);
  signal din1_1_q_net: std_logic_vector(11 downto 0);
  signal din2_0_q_net: std_logic_vector(11 downto 0);
  signal din2_1_q_net: std_logic_vector(11 downto 0);
  signal din2_2_q_net: std_logic_vector(11 downto 0);
  signal din2_3_q_net: std_logic_vector(11 downto 0);
  signal din3_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_2_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_3_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_4_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_5_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_6_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_7_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_8_q_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x35 <= ce_1;
  clk_1_sg_x35 <= clk_1;
  reinterpret1_output_port_net_x3 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_8403f05c85: entity work.bussify_entity_8403f05c85
    port map (
      in1 => din3_0_q_net_x0,
      in2 => din3_1_q_net_x0,
      in3 => din3_2_q_net_x0,
      in4 => din3_3_q_net_x0,
      in5 => din3_4_q_net_x0,
      in6 => din3_5_q_net_x0,
      in7 => din3_6_q_net_x0,
      in8 => din3_7_q_net_x0,
      in9 => din3_8_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => reinterpret1_output_port_net_x3,
      en => '1',
      rst => '1',
      q => din0_0_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_0_q_net
    );

  din1_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_1_q_net
    );

  din2_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din1_0_q_net,
      en => '1',
      rst => '1',
      q => din2_0_q_net
    );

  din2_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din1_1_q_net,
      en => '1',
      rst => '1',
      q => din2_1_q_net
    );

  din2_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din1_0_q_net,
      en => '1',
      rst => '1',
      q => din2_2_q_net
    );

  din2_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din1_1_q_net,
      en => '1',
      rst => '1',
      q => din2_3_q_net
    );

  din3_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_0_q_net,
      en => '1',
      rst => '1',
      q => din3_0_q_net_x0
    );

  din3_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_1_q_net,
      en => '1',
      rst => '1',
      q => din3_1_q_net_x0
    );

  din3_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_2_q_net,
      en => '1',
      rst => '1',
      q => din3_2_q_net_x0
    );

  din3_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_3_q_net,
      en => '1',
      rst => '1',
      q => din3_3_q_net_x0
    );

  din3_4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_0_q_net,
      en => '1',
      rst => '1',
      q => din3_4_q_net_x0
    );

  din3_5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_1_q_net,
      en => '1',
      rst => '1',
      q => din3_5_q_net_x0
    );

  din3_6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_2_q_net,
      en => '1',
      rst => '1',
      q => din3_6_q_net_x0
    );

  din3_7: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_3_q_net,
      en => '1',
      rst => '1',
      q => din3_7_q_net_x0
    );

  din3_8: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      d => din2_0_q_net,
      en => '1',
      rst => '1',
      q => din3_8_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/rep_we/bussify"

entity bussify_entity_66a706537c is
  port (
    in1: in std_logic; 
    in2: in std_logic; 
    in3: in std_logic; 
    in4: in std_logic; 
    in5: in std_logic; 
    in6: in std_logic; 
    in7: in std_logic; 
    in8: in std_logic; 
    in9: in std_logic; 
    bus_out: out std_logic_vector(8 downto 0)
  );
end bussify_entity_66a706537c;

architecture structural of bussify_entity_66a706537c is
  signal concatenate_y_net_x1: std_logic_vector(8 downto 0);
  signal din3_0_q_net_x0: std_logic;
  signal din3_1_q_net_x0: std_logic;
  signal din3_2_q_net_x0: std_logic;
  signal din3_3_q_net_x0: std_logic;
  signal din3_4_q_net_x0: std_logic;
  signal din3_5_q_net_x0: std_logic;
  signal din3_6_q_net_x0: std_logic;
  signal din3_7_q_net_x0: std_logic;
  signal din3_8_q_net_x0: std_logic;
  signal reinterpret1_output_port_net: std_logic;
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic;
  signal reinterpret4_output_port_net: std_logic;
  signal reinterpret5_output_port_net: std_logic;
  signal reinterpret6_output_port_net: std_logic;
  signal reinterpret7_output_port_net: std_logic;
  signal reinterpret8_output_port_net: std_logic;
  signal reinterpret9_output_port_net: std_logic;

begin
  din3_0_q_net_x0 <= in1;
  din3_1_q_net_x0 <= in2;
  din3_2_q_net_x0 <= in3;
  din3_3_q_net_x0 <= in4;
  din3_4_q_net_x0 <= in5;
  din3_5_q_net_x0 <= in6;
  din3_6_q_net_x0 <= in7;
  din3_7_q_net_x0 <= in8;
  din3_8_q_net_x0 <= in9;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_0cc72cd991
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2(0) => reinterpret3_output_port_net,
      in3(0) => reinterpret4_output_port_net,
      in4(0) => reinterpret5_output_port_net,
      in5(0) => reinterpret6_output_port_net,
      in6(0) => reinterpret7_output_port_net,
      in7(0) => reinterpret8_output_port_net,
      in8(0) => reinterpret9_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_0_q_net_x0,
      output_port(0) => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_1_q_net_x0,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_2_q_net_x0,
      output_port(0) => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_3_q_net_x0,
      output_port(0) => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_4_q_net_x0,
      output_port(0) => reinterpret5_output_port_net
    );

  reinterpret6: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_5_q_net_x0,
      output_port(0) => reinterpret6_output_port_net
    );

  reinterpret7: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_6_q_net_x0,
      output_port(0) => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_7_q_net_x0,
      output_port(0) => reinterpret8_output_port_net
    );

  reinterpret9: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_8_q_net_x0,
      output_port(0) => reinterpret9_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0/rep_we"

entity rep_we_entity_e501618f96 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic_vector(8 downto 0)
  );
end rep_we_entity_e501618f96;

architecture structural of rep_we_entity_e501618f96 is
  signal ce_1_sg_x36: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(8 downto 0);
  signal din0_0_q_net: std_logic;
  signal din1_0_q_net: std_logic;
  signal din1_1_q_net: std_logic;
  signal din2_0_q_net: std_logic;
  signal din2_1_q_net: std_logic;
  signal din2_2_q_net: std_logic;
  signal din2_3_q_net: std_logic;
  signal din3_0_q_net_x0: std_logic;
  signal din3_1_q_net_x0: std_logic;
  signal din3_2_q_net_x0: std_logic;
  signal din3_3_q_net_x0: std_logic;
  signal din3_4_q_net_x0: std_logic;
  signal din3_5_q_net_x0: std_logic;
  signal din3_6_q_net_x0: std_logic;
  signal din3_7_q_net_x0: std_logic;
  signal din3_8_q_net_x0: std_logic;
  signal slice1_y_net_x0: std_logic;

begin
  ce_1_sg_x36 <= ce_1;
  clk_1_sg_x36 <= clk_1;
  slice1_y_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_66a706537c: entity work.bussify_entity_66a706537c
    port map (
      in1 => din3_0_q_net_x0,
      in2 => din3_1_q_net_x0,
      in3 => din3_2_q_net_x0,
      in4 => din3_3_q_net_x0,
      in5 => din3_4_q_net_x0,
      in6 => din3_5_q_net_x0,
      in7 => din3_6_q_net_x0,
      in8 => din3_7_q_net_x0,
      in9 => din3_8_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => slice1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_0_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din0_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_0_q_net
    );

  din1_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din0_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_1_q_net
    );

  din2_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din1_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din2_0_q_net
    );

  din2_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din1_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din2_1_q_net
    );

  din2_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din1_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din2_2_q_net
    );

  din2_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din1_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din2_3_q_net
    );

  din3_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_0_q_net_x0
    );

  din3_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_1_q_net_x0
    );

  din3_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_2_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_2_q_net_x0
    );

  din3_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_3_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_3_q_net_x0
    );

  din3_4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_4_q_net_x0
    );

  din3_5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_5_q_net_x0
    );

  din3_6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_2_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_6_q_net_x0
    );

  din3_7: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_3_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_7_q_net_x0
    );

  din3_8: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => din2_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din3_8_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/buf0"

entity buf0_entity_136f881010 is
  port (
    addr: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    we: in std_logic; 
    dout: out std_logic_vector(35 downto 0)
  );
end buf0_entity_136f881010;

architecture structural of buf0_entity_136f881010 is
  signal bram0_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram4_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram5_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram6_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram7_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram8_data_out_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x37: std_logic;
  signal clk_1_sg_x37: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(107 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(8 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(35 downto 0);
  signal ddin_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_din0_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret5_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret5_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret6_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret6_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret7_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret7_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret8_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret8_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret9_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret9_output_port_net_x1: std_logic_vector(3 downto 0);
  signal slice1_y_net_x0: std_logic;
  signal slice1_y_net_x2: std_logic;
  signal slice2_y_net_x0: std_logic;
  signal slice3_y_net_x0: std_logic;
  signal slice4_y_net_x0: std_logic;
  signal slice5_y_net_x0: std_logic;
  signal slice6_y_net_x0: std_logic;
  signal slice7_y_net_x0: std_logic;
  signal slice8_y_net_x0: std_logic;
  signal slice9_y_net_x0: std_logic;

begin
  reinterpret1_output_port_net_x5 <= addr;
  ce_1_sg_x37 <= ce_1;
  clk_1_sg_x37 <= clk_1;
  delay_din0_q_net_x0 <= din;
  slice1_y_net_x2 <= we;
  dout <= concatenate_y_net_x4;

  bram0: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret9_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret9_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice9_y_net_x0,
      data_out => bram0_data_out_net_x0
    );

  bram1: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret8_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret8_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice8_y_net_x0,
      data_out => bram1_data_out_net_x0
    );

  bram2: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret7_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret7_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice7_y_net_x0,
      data_out => bram2_data_out_net_x0
    );

  bram3: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret6_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret6_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice6_y_net_x0,
      data_out => bram3_data_out_net_x0
    );

  bram4: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret5_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret5_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice5_y_net_x0,
      data_out => bram4_data_out_net_x0
    );

  bram5: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret4_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret4_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice4_y_net_x0,
      data_out => bram5_data_out_net_x0
    );

  bram6: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret3_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret3_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice3_y_net_x0,
      data_out => bram6_data_out_net_x0
    );

  bram7: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret2_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret2_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice2_y_net_x0,
      data_out => bram7_data_out_net_x0
    );

  bram8: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      data_in => reinterpret1_output_port_net_x4,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram8_data_out_net_x0
    );

  ddin: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      clr => '0',
      d => delay_din0_q_net_x0,
      q => ddin_q_net_x0
    );

  debus_addr_683e5a971d: entity work.debus_addr_entity_683e5a971d
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out9 => reinterpret9_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0,
      out4 => reinterpret4_output_port_net_x0,
      out5 => reinterpret5_output_port_net_x0,
      out6 => reinterpret6_output_port_net_x0,
      out7 => reinterpret7_output_port_net_x0,
      out8 => reinterpret8_output_port_net_x0
    );

  debus_din_d2fe8dc95c: entity work.debus_din_entity_d2fe8dc95c
    port map (
      bus_in => ddin_q_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out9 => reinterpret9_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1,
      out4 => reinterpret4_output_port_net_x1,
      out5 => reinterpret5_output_port_net_x1,
      out6 => reinterpret6_output_port_net_x1,
      out7 => reinterpret7_output_port_net_x1,
      out8 => reinterpret8_output_port_net_x1
    );

  debus_we_118daa2628: entity work.debus_we_entity_118daa2628
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => slice1_y_net_x0,
      msb_out9 => slice9_y_net_x0,
      out2 => slice2_y_net_x0,
      out3 => slice3_y_net_x0,
      out4 => slice4_y_net_x0,
      out5 => slice5_y_net_x0,
      out6 => slice6_y_net_x0,
      out7 => slice7_y_net_x0,
      out8 => slice8_y_net_x0
    );

  din_bussify_e936a8b4d0: entity work.din_bussify_entity_e936a8b4d0
    port map (
      in1 => bram0_data_out_net_x0,
      in2 => bram1_data_out_net_x0,
      in3 => bram2_data_out_net_x0,
      in4 => bram3_data_out_net_x0,
      in5 => bram4_data_out_net_x0,
      in6 => bram5_data_out_net_x0,
      in7 => bram6_data_out_net_x0,
      in8 => bram7_data_out_net_x0,
      in9 => bram8_data_out_net_x0,
      bus_out => concatenate_y_net_x4
    );

  rep_addr_152c8d6b28: entity work.rep_addr_entity_152c8d6b28
    port map (
      ce_1 => ce_1_sg_x37,
      clk_1 => clk_1_sg_x37,
      in_x0 => reinterpret1_output_port_net_x5,
      out_x0 => concatenate_y_net_x2
    );

  rep_we_e501618f96: entity work.rep_we_entity_e501618f96
    port map (
      ce_1 => ce_1_sg_x37,
      clk_1 => clk_1_sg_x37,
      in_x0 => slice1_y_net_x2,
      out_x0 => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/sync_delay_en"

entity sync_delay_en_entity_5c657e9304 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_en_entity_5c657e9304;

architecture structural of sync_delay_en_entity_5c657e9304 is
  signal ce_1_sg_x38: std_logic;
  signal clk_1_sg_x38: std_logic;
  signal constant1_op_net: std_logic_vector(12 downto 0);
  signal constant2_op_net: std_logic_vector(12 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal logical1_y_net: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x0: std_logic;
  signal or_y_net_x0: std_logic;
  signal pre_sync_delay_q_net_x0: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x38 <= ce_1;
  clk_1_sg_x38 <= clk_1;
  or_y_net_x0 <= en;
  pre_sync_delay_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x0;

  constant1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_50be3b5040
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_eb4d9e2dad
    port map (
      ce => ce_1_sg_x38,
      clk => clk_1_sg_x38,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical1_y_net,
      load(0) => pre_sync_delay_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net,
      d1(0) => or_y_net_x0,
      y(0) => logical1_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x0
    );

  relational: entity work.relational_6dfa374756
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_2550da35d2
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even/we_expand"

entity we_expand_entity_d31ff06e83 is
  port (
    bus_in: in std_logic; 
    msb_lsb_out1: out std_logic
  );
end we_expand_entity_d31ff06e83;

architecture structural of we_expand_entity_d31ff06e83 is
  signal reinterpret1_output_port_net_x0: std_logic;
  signal slice1_y_net_x3: std_logic;

begin
  reinterpret1_output_port_net_x0 <= bus_in;
  msb_lsb_out1 <= slice1_y_net_x3;

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 1,
      y_width => 1
    )
    port map (
      x(0) => reinterpret1_output_port_net_x0,
      y(0) => slice1_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_even"

entity reorder_even_entity_db2ff2e020 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end reorder_even_entity_db2ff2e020;

architecture structural of reorder_even_entity_db2ff2e020 is
  signal ce_1_sg_x39: std_logic;
  signal clk_1_sg_x39: std_logic;
  signal concatenate_y_net_x5: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we0_q_net: std_logic;
  signal delay_we2_q_net_x1: std_logic;
  signal en_even_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic;
  signal mux_y_net_x1: std_logic_vector(11 downto 0);
  signal or_y_net_x0: std_logic;
  signal post_sync_delay_q_net_x0: std_logic;
  signal pre_sync_delay_q_net_x0: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic;
  signal reinterpret1_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice1_y_net_x3: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x39 <= ce_1;
  clk_1_sg_x39 <= clk_1;
  reinterpret2_output_port_net_x0 <= din0;
  en_even_op_net_x0 <= en;
  delay0_q_net_x0 <= sync;
  dout0 <= concatenate_y_net_x5;
  sync_out <= post_sync_delay_q_net_x0;

  addr_expand_8d8c5a295c: entity work.addr_expand_entity_8d8c5a295c
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x5
    );

  addr_replicate_cc9047aff8: entity work.addr_replicate_entity_cc9047aff8
    port map (
      in_x0 => mux_y_net_x1,
      out_x0 => reinterpret1_output_port_net_x3
    );

  buf0_136f881010: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret1_output_port_net_x5,
      ce_1 => ce_1_sg_x39,
      clk_1 => clk_1_sg_x39,
      din => delay_din0_q_net_x0,
      we => slice1_y_net_x3,
      dout => concatenate_y_net_x5
    );

  counter: entity work.counter_486acbf0b9
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      en(0) => en_even_op_net_x0,
      rst(0) => delay0_q_net_x0,
      op => counter_op_net
    );

  delay_d0: entity work.delay_b1290993d1
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d => reinterpret2_output_port_net_x0,
      q => delay_din0_q_net_x0
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_85c2ef968b
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we0: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d(0) => en_even_op_net_x0,
      q(0) => delay_we0_q_net
    );

  delay_we2: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d(0) => en_even_op_net_x0,
      q(0) => delay_we2_q_net_x1
    );

  map1: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 12,
      core_name0 => "bmg_72_180432cd81ea5a8d",
      latency => 2
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      en => "1",
      rst => "0",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net_x1
    );

  or_x0: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => pre_sync_delay_q_net_x0,
      d1(0) => delay_we0_q_net,
      y(0) => or_y_net_x0
    );

  post_sync_delay: entity work.delay_fa260f7d22
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => post_sync_delay_q_net_x0
    );

  pre_sync_delay: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      clr => '0',
      d(0) => delay0_q_net_x0,
      q(0) => pre_sync_delay_q_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

  sync_delay_en_5c657e9304: entity work.sync_delay_en_entity_5c657e9304
    port map (
      ce_1 => ce_1_sg_x39,
      clk_1 => clk_1_sg_x39,
      en => or_y_net_x0,
      in_x0 => pre_sync_delay_q_net_x0,
      out_x0 => mux_y_net_x0
    );

  we_expand_d31ff06e83: entity work.we_expand_entity_d31ff06e83
    port map (
      bus_in => reinterpret1_output_port_net_x2,
      msb_lsb_out1 => slice1_y_net_x3
    );

  we_replicate_63f30adcba: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => delay_we2_q_net_x1,
      out_x0 => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_odd"

entity reorder_odd_entity_e91138e8d9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0)
  );
end reorder_odd_entity_e91138e8d9;

architecture structural of reorder_odd_entity_e91138e8d9 is
  signal ce_1_sg_x43: std_logic;
  signal clk_1_sg_x43: std_logic;
  signal concatenate_y_net_x5: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we2_q_net_x1: std_logic;
  signal en_odd_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net_x1: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic;
  signal reinterpret1_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(11 downto 0);
  signal slice1_y_net: std_logic;
  signal slice1_y_net_x3: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x43 <= ce_1;
  clk_1_sg_x43 <= clk_1;
  reinterpret1_output_port_net_x0 <= din0;
  en_odd_op_net_x0 <= en;
  delay0_q_net_x1 <= sync;
  dout0 <= concatenate_y_net_x5;

  addr_expand_a4272c8866: entity work.addr_expand_entity_8d8c5a295c
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x5
    );

  addr_replicate_f5d7bc66c1: entity work.addr_replicate_entity_cc9047aff8
    port map (
      in_x0 => mux_y_net_x1,
      out_x0 => reinterpret1_output_port_net_x3
    );

  buf0_3524aa9016: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret1_output_port_net_x5,
      ce_1 => ce_1_sg_x43,
      clk_1 => clk_1_sg_x43,
      din => delay_din0_q_net_x0,
      we => slice1_y_net_x3,
      dout => concatenate_y_net_x5
    );

  counter: entity work.counter_486acbf0b9
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      en(0) => en_odd_op_net_x0,
      rst(0) => delay0_q_net_x1,
      op => counter_op_net
    );

  delay_d0: entity work.delay_b1290993d1
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => delay_din0_q_net_x0
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_85c2ef968b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we2: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      d(0) => en_odd_op_net_x0,
      q(0) => delay_we2_q_net_x1
    );

  map1: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 12,
      core_name0 => "bmg_72_8574240a262aac9a",
      latency => 2
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      en => "1",
      rst => "0",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

  we_expand_743d567645: entity work.we_expand_entity_d31ff06e83
    port map (
      bus_in => reinterpret1_output_port_net_x2,
      msb_lsb_out1 => slice1_y_net_x3
    );

  we_replicate_17836f8c07: entity work.sel_replicate0_entity_bc92d7dfef
    port map (
      in_x0 => delay_we2_q_net_x1,
      out_x0 => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/addr_expand"

entity addr_expand_entity_80b50b7dd2 is
  port (
    bus_in: in std_logic_vector(47 downto 0); 
    lsb_out1: out std_logic_vector(11 downto 0); 
    msb_out4: out std_logic_vector(11 downto 0); 
    out2: out std_logic_vector(11 downto 0); 
    out3: out std_logic_vector(11 downto 0)
  );
end addr_expand_entity_80b50b7dd2;

architecture structural of addr_expand_entity_80b50b7dd2 is
  signal concatenate_y_net_x0: std_logic_vector(47 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(11 downto 0);
  signal slice1_y_net: std_logic_vector(11 downto 0);
  signal slice2_y_net: std_logic_vector(11 downto 0);
  signal slice3_y_net: std_logic_vector(11 downto 0);
  signal slice4_y_net: std_logic_vector(11 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 48,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 23,
      x_width => 48,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 35,
      x_width => 48,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 47,
      x_width => 48,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/addr_replicate/bussify"

entity bussify_entity_d7ecf11fe9 is
  port (
    in1: in std_logic_vector(11 downto 0); 
    in2: in std_logic_vector(11 downto 0); 
    in3: in std_logic_vector(11 downto 0); 
    in4: in std_logic_vector(11 downto 0); 
    bus_out: out std_logic_vector(47 downto 0)
  );
end bussify_entity_d7ecf11fe9;

architecture structural of bussify_entity_d7ecf11fe9 is
  signal concatenate_y_net_x1: std_logic_vector(47 downto 0);
  signal din1_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_2_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_3_q_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(11 downto 0);

begin
  din1_0_q_net_x0 <= in1;
  din1_1_q_net_x0 <= in2;
  din1_2_q_net_x0 <= in3;
  din1_3_q_net_x0 <= in4;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_08ed6107eb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din1_0_q_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din1_1_q_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din1_2_q_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din1_3_q_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/addr_replicate"

entity addr_replicate_entity_d68dbd7454 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(47 downto 0)
  );
end addr_replicate_entity_d68dbd7454;

architecture structural of addr_replicate_entity_d68dbd7454 is
  signal ce_1_sg_x44: std_logic;
  signal clk_1_sg_x44: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(47 downto 0);
  signal din0_0_q_net: std_logic_vector(11 downto 0);
  signal din0_1_q_net: std_logic_vector(11 downto 0);
  signal din1_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_2_q_net_x0: std_logic_vector(11 downto 0);
  signal din1_3_q_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x44 <= ce_1;
  clk_1_sg_x44 <= clk_1;
  mux_y_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_d7ecf11fe9: entity work.bussify_entity_d7ecf11fe9
    port map (
      in1 => din1_0_q_net_x0,
      in2 => din1_1_q_net_x0,
      in3 => din1_2_q_net_x0,
      in4 => din1_3_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => mux_y_net_x0,
      en => '1',
      rst => '1',
      q => din0_0_q_net
    );

  din0_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => mux_y_net_x0,
      en => '1',
      rst => '1',
      q => din0_1_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_0_q_net_x0
    );

  din1_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => din0_1_q_net,
      en => '1',
      rst => '1',
      q => din1_1_q_net_x0
    );

  din1_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_2_q_net_x0
    );

  din1_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      d => din0_1_q_net,
      en => '1',
      rst => '1',
      q => din1_3_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/we_expand"

entity we_expand_entity_89eef2f68f is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    lsb_out1: out std_logic; 
    msb_out4: out std_logic; 
    out2: out std_logic; 
    out3: out std_logic
  );
end we_expand_entity_89eef2f68f;

architecture structural of we_expand_entity_89eef2f68f is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net_x3: std_logic;
  signal slice2_y_net_x3: std_logic;
  signal slice3_y_net_x3: std_logic;
  signal slice4_y_net_x3: std_logic;

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= slice1_y_net_x3;
  msb_out4 <= slice4_y_net_x3;
  out2 <= slice2_y_net_x3;
  out3 <= slice3_y_net_x3;

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice1_y_net_x3
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice2_y_net_x3
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice3_y_net_x3
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice4_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/we_replicate/bussify"

entity bussify_entity_6bd38bcd1d is
  port (
    in1: in std_logic; 
    in2: in std_logic; 
    in3: in std_logic; 
    in4: in std_logic; 
    bus_out: out std_logic_vector(3 downto 0)
  );
end bussify_entity_6bd38bcd1d;

architecture structural of bussify_entity_6bd38bcd1d is
  signal concatenate_y_net_x1: std_logic_vector(3 downto 0);
  signal din1_0_q_net_x0: std_logic;
  signal din1_1_q_net_x0: std_logic;
  signal din1_2_q_net_x0: std_logic;
  signal din1_3_q_net_x0: std_logic;
  signal reinterpret1_output_port_net: std_logic;
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic;
  signal reinterpret4_output_port_net: std_logic;

begin
  din1_0_q_net_x0 <= in1;
  din1_1_q_net_x0 <= in2;
  din1_2_q_net_x0 <= in3;
  din1_3_q_net_x0 <= in4;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2(0) => reinterpret3_output_port_net,
      in3(0) => reinterpret4_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din1_0_q_net_x0,
      output_port(0) => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din1_1_q_net_x0,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din1_2_q_net_x0,
      output_port(0) => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din1_3_q_net_x0,
      output_port(0) => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out/we_replicate"

entity we_replicate_entity_35844a72d5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic_vector(3 downto 0)
  );
end we_replicate_entity_35844a72d5;

architecture structural of we_replicate_entity_35844a72d5 is
  signal ce_1_sg_x57: std_logic;
  signal clk_1_sg_x57: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(3 downto 0);
  signal delay_we2_q_net_x0: std_logic;
  signal din0_0_q_net: std_logic;
  signal din0_1_q_net: std_logic;
  signal din1_0_q_net_x0: std_logic;
  signal din1_1_q_net_x0: std_logic;
  signal din1_2_q_net_x0: std_logic;
  signal din1_3_q_net_x0: std_logic;

begin
  ce_1_sg_x57 <= ce_1;
  clk_1_sg_x57 <= clk_1;
  delay_we2_q_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_6bd38bcd1d: entity work.bussify_entity_6bd38bcd1d
    port map (
      in1 => din1_0_q_net_x0,
      in2 => din1_1_q_net_x0,
      in3 => din1_2_q_net_x0,
      in4 => din1_3_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => delay_we2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_0_q_net
    );

  din0_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => delay_we2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_1_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => din0_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_0_q_net_x0
    );

  din1_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => din0_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_1_q_net_x0
    );

  din1_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => din0_0_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_2_q_net_x0
    );

  din1_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => din0_1_q_net,
      en => '1',
      rst => '1',
      q(0) => din1_3_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/reorder_out"

entity reorder_out_entity_22c6aa5a0c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din0: in std_logic_vector(35 downto 0); 
    din1: in std_logic_vector(35 downto 0); 
    din2: in std_logic_vector(35 downto 0); 
    din3: in std_logic_vector(35 downto 0); 
    en: in std_logic; 
    sync: in std_logic; 
    dout0: out std_logic_vector(35 downto 0); 
    dout1: out std_logic_vector(35 downto 0); 
    dout2: out std_logic_vector(35 downto 0); 
    dout3: out std_logic_vector(35 downto 0)
  );
end reorder_out_entity_22c6aa5a0c;

architecture structural of reorder_out_entity_22c6aa5a0c is
  signal ce_1_sg_x58: std_logic;
  signal clk_1_sg_x58: std_logic;
  signal concatenate_y_net_x10: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(47 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay_d0_q_net: std_logic_vector(11 downto 0);
  signal delay_din0_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_din1_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_din2_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_din3_q_net_x0: std_logic_vector(35 downto 0);
  signal delay_map1_q_net: std_logic_vector(11 downto 0);
  signal delay_sel_q_net: std_logic;
  signal delay_we2_q_net_x0: std_logic;
  signal en_out_op_net_x0: std_logic;
  signal map1_data_net: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x2: std_logic;
  signal ram_data_out_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret4_output_port_net_x3: std_logic_vector(11 downto 0);
  signal reinterpret_out_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x13: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic;
  signal slice1_y_net_x3: std_logic;
  signal slice2_y_net: std_logic_vector(11 downto 0);
  signal slice2_y_net_x3: std_logic;
  signal slice3_y_net_x3: std_logic;
  signal slice4_y_net_x3: std_logic;

begin
  ce_1_sg_x58 <= ce_1;
  clk_1_sg_x58 <= clk_1;
  ram_data_out_net_x4 <= din0;
  ram_data_out_net_x5 <= din1;
  reinterpret_out_output_port_net_x12 <= din2;
  reinterpret_out_output_port_net_x13 <= din3;
  en_out_op_net_x0 <= en;
  mux_y_net_x2 <= sync;
  dout0 <= concatenate_y_net_x9;
  dout1 <= concatenate_y_net_x10;
  dout2 <= concatenate_y_net_x11;
  dout3 <= concatenate_y_net_x12;

  addr_expand_80b50b7dd2: entity work.addr_expand_entity_80b50b7dd2
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x3,
      msb_out4 => reinterpret4_output_port_net_x3,
      out2 => reinterpret2_output_port_net_x3,
      out3 => reinterpret3_output_port_net_x3
    );

  addr_replicate_d68dbd7454: entity work.addr_replicate_entity_d68dbd7454
    port map (
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      in_x0 => mux_y_net_x0,
      out_x0 => concatenate_y_net_x2
    );

  buf0_896c373683: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret4_output_port_net_x3,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => delay_din0_q_net_x0,
      we => slice4_y_net_x3,
      dout => concatenate_y_net_x9
    );

  buf1_8ea2217a94: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret3_output_port_net_x3,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => delay_din1_q_net_x0,
      we => slice3_y_net_x3,
      dout => concatenate_y_net_x10
    );

  buf2_6d8ff8cf4d: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => delay_din2_q_net_x0,
      we => slice2_y_net_x3,
      dout => concatenate_y_net_x11
    );

  buf3_d026baa734: entity work.buf0_entity_136f881010
    port map (
      addr => reinterpret1_output_port_net_x3,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      din => delay_din3_q_net_x0,
      we => slice1_y_net_x3,
      dout => concatenate_y_net_x12
    );

  counter: entity work.counter_486acbf0b9
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      en(0) => en_out_op_net_x0,
      rst(0) => mux_y_net_x2,
      op => counter_op_net
    );

  delay_d0: entity work.delay_b1290993d1
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d => slice2_y_net,
      q => delay_d0_q_net
    );

  delay_din0: entity work.delay_28d2c9d50c
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d => ram_data_out_net_x4,
      q => delay_din0_q_net_x0
    );

  delay_din1: entity work.delay_28d2c9d50c
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d => ram_data_out_net_x5,
      q => delay_din1_q_net_x0
    );

  delay_din2: entity work.delay_28d2c9d50c
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d => reinterpret_out_output_port_net_x12,
      q => delay_din2_q_net_x0
    );

  delay_din3: entity work.delay_28d2c9d50c
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d => reinterpret_out_output_port_net_x13,
      q => delay_din3_q_net_x0
    );

  delay_map1: entity work.delay_4670f4967f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => map1_data_net,
      q => delay_map1_q_net
    );

  delay_sel: entity work.delay_85c2ef968b
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d(0) => slice1_y_net,
      q(0) => delay_sel_q_net
    );

  delay_we2: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d(0) => en_out_op_net_x0,
      q(0) => delay_we2_q_net_x0
    );

  map1: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 12,
      core_name0 => "bmg_72_ce7e9961dfcc2802",
      latency => 2
    )
    port map (
      addr => slice2_y_net,
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      en => "1",
      rst => "0",
      data => map1_data_net
    );

  mux: entity work.mux_25f2d74a2a
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      d0 => delay_d0_q_net,
      d1 => delay_map1_q_net,
      sel(0) => delay_sel_q_net,
      y => mux_y_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 13,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice2_y_net
    );

  we_expand_89eef2f68f: entity work.we_expand_entity_89eef2f68f
    port map (
      bus_in => concatenate_y_net_x8,
      lsb_out1 => slice1_y_net_x3,
      msb_out4 => slice4_y_net_x3,
      out2 => slice2_y_net_x3,
      out3 => slice3_y_net_x3
    );

  we_replicate_35844a72d5: entity work.we_replicate_entity_35844a72d5
    port map (
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      in_x0 => delay_we2_q_net_x0,
      out_x0 => concatenate_y_net_x8
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x/sync_delay"

entity sync_delay_entity_c43fa8c0d9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_c43fa8c0d9;

architecture structural of sync_delay_entity_c43fa8c0d9 is
  signal ce_1_sg_x59: std_logic;
  signal clk_1_sg_x59: std_logic;
  signal constant1_op_net: std_logic_vector(12 downto 0);
  signal constant2_op_net: std_logic_vector(12 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(12 downto 0);
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal d2_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x3: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x59 <= ce_1;
  clk_1_sg_x59 <= clk_1;
  d2_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x3;

  constant1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_50be3b5040
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_eb4d9e2dad
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => d2_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => d2_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => d2_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x3
    );

  relational: entity work.relational_6dfa374756
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_2550da35d2
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/bi_real_unscr_4x"

entity bi_real_unscr_4x_entity_b9d413eca4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    even: in std_logic_vector(35 downto 0); 
    odd: in std_logic_vector(35 downto 0); 
    sync: in std_logic; 
    pol1_out: out std_logic_vector(35 downto 0); 
    pol2_out: out std_logic_vector(35 downto 0); 
    pol3_out: out std_logic_vector(35 downto 0); 
    pol4_out: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end bi_real_unscr_4x_entity_b9d413eca4;

architecture structural of bi_real_unscr_4x_entity_b9d413eca4 is
  signal c0_op_net: std_logic_vector(12 downto 0);
  signal c1_op_net: std_logic_vector(12 downto 0);
  signal ce_1_sg_x60: std_logic;
  signal clk_1_sg_x60: std_logic;
  signal concatenate_y_net_x10: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(35 downto 0);
  signal count_op_net: std_logic_vector(12 downto 0);
  signal d0_q_net: std_logic_vector(35 downto 0);
  signal d2_q_net_x0: std_logic;
  signal d3_q_net_x2: std_logic_vector(35 downto 0);
  signal d4_q_net_x2: std_logic_vector(35 downto 0);
  signal d5_q_net_x2: std_logic_vector(35 downto 0);
  signal d6_q_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal en_even_op_net_x0: std_logic;
  signal en_odd_op_net_x0: std_logic;
  signal en_out_op_net_x0: std_logic;
  signal mux0_y_net_x1: std_logic_vector(35 downto 0);
  signal mux1_y_net_x1: std_logic_vector(35 downto 0);
  signal mux2_y_net_x1: std_logic_vector(35 downto 0);
  signal mux3_y_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal post_sync_delay_q_net_x0: std_logic;
  signal r0_op_net: std_logic;
  signal r1_op_net: std_logic;
  signal ram_data_out_net_x4: std_logic_vector(35 downto 0);
  signal ram_data_out_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x18: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x19: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x20: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x21: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x22: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x13: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x6: std_logic_vector(35 downto 0);
  signal sync_delay1_q_net_x1: std_logic;

begin
  ce_1_sg_x60 <= ce_1;
  clk_1_sg_x60 <= clk_1;
  reinterpret2_output_port_net_x1 <= even;
  reinterpret1_output_port_net_x18 <= odd;
  delay0_q_net_x2 <= sync;
  pol1_out <= reinterpret1_output_port_net_x19;
  pol2_out <= reinterpret1_output_port_net_x20;
  pol3_out <= reinterpret1_output_port_net_x21;
  pol4_out <= reinterpret1_output_port_net_x22;
  sync_out <= sync_delay1_q_net_x1;

  c0: entity work.constant_e47f8076b8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => c0_op_net
    );

  c1: entity work.constant_0c8736a503
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => c1_op_net
    );

  count: entity work.counter_c48d6dcab5
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      rst(0) => post_sync_delay_q_net_x0,
      op => count_op_net
    );

  d0: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d => concatenate_y_net_x6,
      q => d0_q_net
    );

  d2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d(0) => post_sync_delay_q_net_x0,
      q(0) => d2_q_net_x0
    );

  d3: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d => concatenate_y_net_x9,
      q => d3_q_net_x2
    );

  d4: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d => concatenate_y_net_x10,
      q => d4_q_net_x2
    );

  d5: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d => concatenate_y_net_x11,
      q => d5_q_net_x2
    );

  d6: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d => concatenate_y_net_x12,
      q => d6_q_net_x2
    );

  delay0_f75f886771: entity work.delay0_entity_f75f886771
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din => reinterpret_out_output_port_net_x5,
      dout => ram_data_out_net_x4
    );

  delay1_0843e4dc11: entity work.delay0_entity_f75f886771
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din => reinterpret_out_output_port_net_x6,
      dout => ram_data_out_net_x5
    );

  en_even: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_even_op_net_x0
    );

  en_odd: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_odd_op_net_x0
    );

  en_out: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => en_out_op_net_x0
    );

  hilbert0_99acf82149: entity work.hilbert0_entity_99acf82149
    port map (
      a => mux0_y_net_x1,
      b => mux1_y_net_x1,
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      even => reinterpret_out_output_port_net_x5,
      odd => reinterpret_out_output_port_net_x6
    );

  hilbert1_9cb7ed5b0e: entity work.hilbert0_entity_99acf82149
    port map (
      a => mux2_y_net_x1,
      b => mux3_y_net_x1,
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      even => reinterpret_out_output_port_net_x12,
      odd => reinterpret_out_output_port_net_x13
    );

  mirror_spectrum_dc7f261b12: entity work.mirror_spectrum_entity_dc7f261b12
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din0 => ram_data_out_net_x4,
      din1 => ram_data_out_net_x5,
      din2 => reinterpret_out_output_port_net_x12,
      din3 => reinterpret_out_output_port_net_x13,
      reo_in0 => d3_q_net_x2,
      reo_in1 => d4_q_net_x2,
      reo_in2 => d5_q_net_x2,
      reo_in3 => d6_q_net_x2,
      sync => mux_y_net_x3,
      dout0 => reinterpret1_output_port_net_x19,
      dout1 => reinterpret1_output_port_net_x20,
      dout2 => reinterpret1_output_port_net_x21,
      dout3 => reinterpret1_output_port_net_x22,
      sync_out => sync_delay1_q_net_x1
    );

  mux0: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d0 => concatenate_y_net_x5,
      d1 => d0_q_net,
      sel(0) => r0_op_net,
      y => mux0_y_net_x1
    );

  mux1: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d0 => d0_q_net,
      d1 => concatenate_y_net_x5,
      sel(0) => r1_op_net,
      y => mux1_y_net_x1
    );

  mux2: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d0 => concatenate_y_net_x5,
      d1 => d0_q_net,
      sel(0) => r1_op_net,
      y => mux2_y_net_x1
    );

  mux3: entity work.mux_fca786f2ff
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      d0 => d0_q_net,
      d1 => concatenate_y_net_x5,
      sel(0) => r0_op_net,
      y => mux3_y_net_x1
    );

  r0: entity work.relational_6dfa374756
    port map (
      a => c0_op_net,
      b => count_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => r0_op_net
    );

  r1: entity work.relational_6dfa374756
    port map (
      a => count_op_net,
      b => c1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => r1_op_net
    );

  reorder_even_db2ff2e020: entity work.reorder_even_entity_db2ff2e020
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din0 => reinterpret2_output_port_net_x1,
      en => en_even_op_net_x0,
      sync => delay0_q_net_x2,
      dout0 => concatenate_y_net_x5,
      sync_out => post_sync_delay_q_net_x0
    );

  reorder_odd_e91138e8d9: entity work.reorder_odd_entity_e91138e8d9
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din0 => reinterpret1_output_port_net_x18,
      en => en_odd_op_net_x0,
      sync => delay0_q_net_x2,
      dout0 => concatenate_y_net_x6
    );

  reorder_out_22c6aa5a0c: entity work.reorder_out_entity_22c6aa5a0c
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      din0 => ram_data_out_net_x4,
      din1 => ram_data_out_net_x5,
      din2 => reinterpret_out_output_port_net_x12,
      din3 => reinterpret_out_output_port_net_x13,
      en => en_out_op_net_x0,
      sync => mux_y_net_x3,
      dout0 => concatenate_y_net_x9,
      dout1 => concatenate_y_net_x10,
      dout2 => concatenate_y_net_x11,
      dout3 => concatenate_y_net_x12
    );

  sync_delay_c43fa8c0d9: entity work.sync_delay_entity_c43fa8c0d9
    port map (
      ce_1 => ce_1_sg_x60,
      clk_1 => clk_1_sg_x60,
      in_x0 => d2_q_net_x0,
      out_x0 => mux_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_add/a_debus"

entity a_debus_entity_e8ca01a28d is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out2: out std_logic_vector(17 downto 0)
  );
end a_debus_entity_e8ca01a28d;

architecture structural of a_debus_entity_e8ca01a28d is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_add/op_bussify"

entity op_bussify_entity_a6d4bedd3c is
  port (
    in1: in std_logic_vector(18 downto 0); 
    in2: in std_logic_vector(18 downto 0); 
    bus_out: out std_logic_vector(37 downto 0)
  );
end op_bussify_entity_a6d4bedd3c;

architecture structural of op_bussify_entity_a6d4bedd3c is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(37 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(18 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  addsub2_s_net_x0 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_5a12f8f9be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub2_s_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_add"

entity bus_add_entity_a60c7dc670 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(37 downto 0)
  );
end bus_add_entity_a60c7dc670;

architecture structural of bus_add_entity_a60c7dc670 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x61: std_logic;
  signal clk_1_sg_x61: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(37 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x2 <= a;
  dmux0_q_net_x1 <= b;
  ce_1_sg_x61 <= ce_1;
  clk_1_sg_x61 <= clk_1;
  dout <= concatenate_y_net_x3;

  a_debus_e8ca01a28d: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_0b9daa5d24360c6e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_0b9daa5d24360c6e",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_2aade9f6e8: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => dmux0_q_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_a6d4bedd3c: entity work.op_bussify_entity_a6d4bedd3c
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_convert/conv1/convert"

entity convert_entity_0000fb9a02 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(19 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end convert_entity_0000fb9a02;

architecture structural of convert_entity_0000fb9a02 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x62: std_logic;
  signal clk_1_sg_x62: std_logic;
  signal concat_y_net: std_logic_vector(20 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(20 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(19 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x62 <= ce_1;
  clk_1_sg_x62 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 19,
      a_width => 21,
      b_arith => xlUnsigned,
      b_bin_pt => 19,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 22,
      core_name0 => "addsb_11_0_80a4fb0fcb4866f6",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 22,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 18
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x62,
      clk => clk_1_sg_x62,
      clr => '0',
      en => "1",
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_c615d93998
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_convert/conv1"

entity conv1_entity_fdd5d602ff is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(19 downto 0); 
    dout: out std_logic_vector(17 downto 0); 
    of_x0: out std_logic
  );
end conv1_entity_fdd5d602ff;

architecture structural of conv1_entity_fdd5d602ff is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal all_0s_y_net: std_logic;
  signal all_1s_y_net: std_logic;
  signal and_y_net_x0: std_logic;
  signal ce_1_sg_x63: std_logic;
  signal clk_1_sg_x63: std_logic;
  signal invert1_op_net: std_logic;
  signal invert2_op_net: std_logic;
  signal reinterpret4_output_port_net_x1: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic;

begin
  ce_1_sg_x63 <= ce_1;
  clk_1_sg_x63 <= clk_1;
  reinterpret4_output_port_net_x1 <= din;
  dout <= adder_s_net_x5;
  of_x0 <= and_y_net_x0;

  all_0s: entity work.logical_89dc141487
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      d0(0) => invert1_op_net,
      d1(0) => invert2_op_net,
      y(0) => all_0s_y_net
    );

  all_1s: entity work.logical_89dc141487
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      d0(0) => slice1_y_net,
      d1(0) => slice2_y_net,
      y(0) => all_1s_y_net
    );

  and_x0: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => all_0s_y_net,
      d1(0) => all_1s_y_net,
      y(0) => and_y_net_x0
    );

  convert_0000fb9a02: entity work.convert_entity_0000fb9a02
    port map (
      ce_1 => ce_1_sg_x63,
      clk_1 => clk_1_sg_x63,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  invert1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      ip(0) => slice1_y_net,
      op(0) => invert1_op_net
    );

  invert2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      ip(0) => slice2_y_net,
      op(0) => invert2_op_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 19,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 18,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_convert/debus"

entity debus_entity_5abef6bede is
  port (
    bus_in: in std_logic_vector(79 downto 0); 
    lsb_out1: out std_logic_vector(19 downto 0); 
    msb_out4: out std_logic_vector(19 downto 0); 
    out2: out std_logic_vector(19 downto 0); 
    out3: out std_logic_vector(19 downto 0)
  );
end debus_entity_5abef6bede;

architecture structural of debus_entity_5abef6bede is
  signal concatenate_y_net_x0: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic_vector(19 downto 0);
  signal slice2_y_net: std_logic_vector(19 downto 0);
  signal slice3_y_net: std_logic_vector(19 downto 0);
  signal slice4_y_net: std_logic_vector(19 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out4 <= reinterpret4_output_port_net_x2;
  out2 <= reinterpret2_output_port_net_x2;
  out3 <= reinterpret3_output_port_net_x2;

  reinterpret1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  reinterpret3: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x2
    );

  reinterpret4: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 19,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 39,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 59,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 79,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_convert"

entity bus_convert_entity_7b742cca79 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(71 downto 0); 
    overflow: out std_logic_vector(3 downto 0)
  );
end bus_convert_entity_7b742cca79;

architecture structural of bus_convert_entity_7b742cca79 is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal adder_s_net_x8: std_logic_vector(17 downto 0);
  signal and_y_net_x4: std_logic;
  signal and_y_net_x5: std_logic;
  signal and_y_net_x6: std_logic;
  signal and_y_net_x7: std_logic;
  signal ce_1_sg_x70: std_logic;
  signal clk_1_sg_x70: std_logic;
  signal concatenate_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x70 <= ce_1;
  clk_1_sg_x70 <= clk_1;
  concatenate_y_net_x3 <= din;
  dout <= concatenate_y_net_x4;
  overflow <= concatenate_y_net_x5;

  bussify_c46cecb5e4: entity work.bussify_entity_904656ce6f
    port map (
      in1 => adder_s_net_x5,
      in2 => adder_s_net_x6,
      in3 => adder_s_net_x7,
      in4 => adder_s_net_x8,
      bus_out => concatenate_y_net_x4
    );

  conv1_fdd5d602ff: entity work.conv1_entity_fdd5d602ff
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      din => reinterpret4_output_port_net_x2,
      dout => adder_s_net_x5,
      of_x0 => and_y_net_x4
    );

  conv2_66a0616fea: entity work.conv1_entity_fdd5d602ff
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      din => reinterpret3_output_port_net_x2,
      dout => adder_s_net_x6,
      of_x0 => and_y_net_x5
    );

  conv3_9091c89c5b: entity work.conv1_entity_fdd5d602ff
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      din => reinterpret2_output_port_net_x2,
      dout => adder_s_net_x7,
      of_x0 => and_y_net_x6
    );

  conv4_fbf770d51c: entity work.conv1_entity_fdd5d602ff
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      din => reinterpret1_output_port_net_x2,
      dout => adder_s_net_x8,
      of_x0 => and_y_net_x7
    );

  debus_5abef6bede: entity work.debus_entity_5abef6bede
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

  of_bussify_eabf114a17: entity work.bussify_entity_6bd38bcd1d
    port map (
      in1 => and_y_net_x4,
      in2 => and_y_net_x5,
      in3 => and_y_net_x6,
      in4 => and_y_net_x7,
      bus_out => concatenate_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_expand"

entity bus_expand_entity_f69635d38b is
  port (
    bus_in: in std_logic_vector(71 downto 0); 
    lsb_out1: out std_logic_vector(35 downto 0); 
    msb_out2: out std_logic_vector(35 downto 0)
  );
end bus_expand_entity_f69635d38b;

architecture structural of bus_expand_entity_f69635d38b is
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);
  signal slice2_y_net: std_logic_vector(35 downto 0);

begin
  concatenate_y_net_x5 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 72,
      y_width => 36
    )
    port map (
      x => concatenate_y_net_x5,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 71,
      x_width => 72,
      y_width => 36
    )
    port map (
      x => concatenate_y_net_x5,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_norm0/bussify"

entity bussify_entity_c32f93b775 is
  port (
    in1: in std_logic_vector(19 downto 0); 
    in2: in std_logic_vector(19 downto 0); 
    in3: in std_logic_vector(19 downto 0); 
    in4: in std_logic_vector(19 downto 0); 
    bus_out: out std_logic_vector(79 downto 0)
  );
end bussify_entity_c32f93b775;

architecture structural of bussify_entity_c32f93b775 is
  signal concatenate_y_net_x0: std_logic_vector(79 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(19 downto 0);

begin
  conv1_dout_net_x0 <= in1;
  conv2_dout_net_x0 <= in2;
  conv3_dout_net_x0 <= in3;
  conv4_dout_net_x0 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_f86ebb6084
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv1_dout_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv2_dout_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv3_dout_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv4_dout_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_norm0"

entity bus_norm0_entity_74bb60a7d0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_norm0_entity_74bb60a7d0;

architecture structural of bus_norm0_entity_74bb60a7d0 is
  signal ce_1_sg_x71: std_logic;
  signal clk_1_sg_x71: std_logic;
  signal concat_y_net_x1: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(79 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(19 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x71 <= ce_1;
  clk_1_sg_x71 <= clk_1;
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x1;

  bussify_c32f93b775: entity work.bussify_entity_c32f93b775
    port map (
      in1 => conv1_dout_net_x0,
      in2 => conv2_dout_net_x0,
      in3 => conv3_dout_net_x0,
      in4 => conv4_dout_net_x0,
      bus_out => concatenate_y_net_x1
    );

  conv1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din => reinterpret4_output_port_net_x0,
      en => "1",
      dout => conv1_dout_net_x0
    );

  conv2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din => reinterpret3_output_port_net_x0,
      en => "1",
      dout => conv2_dout_net_x0
    );

  conv3: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din => reinterpret2_output_port_net_x0,
      en => "1",
      dout => conv3_dout_net_x0
    );

  conv4: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 19,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 20,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din => reinterpret1_output_port_net_x0,
      en => "1",
      dout => conv4_dout_net_x0
    );

  debus_baf1625fc6: entity work.debus_entity_b713d0483e
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_norm1/conv1"

entity conv1_entity_254c41df9c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(18 downto 0); 
    out_x0: out std_logic_vector(19 downto 0)
  );
end conv1_entity_254c41df9c;

architecture structural of conv1_entity_254c41df9c is
  signal adder_s_net_x4: std_logic_vector(19 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x72: std_logic;
  signal clk_1_sg_x72: std_logic;
  signal concat_y_net: std_logic_vector(19 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(19 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(18 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x72 <= ce_1;
  clk_1_sg_x72 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 19,
      a_width => 20,
      b_arith => xlUnsigned,
      b_bin_pt => 19,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 21,
      core_name0 => "addsb_11_0_3af1276811d12ede",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 21,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 18,
      s_width => 20
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x72,
      clk => clk_1_sg_x72,
      clr => '0',
      en => "1",
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_b366689086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 19,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_504cae28bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_bc4405cd1e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_b1e9d7c303
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_norm1"

entity bus_norm1_entity_b00e4bc012 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(75 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_norm1_entity_b00e4bc012;

architecture structural of bus_norm1_entity_b00e4bc012 is
  signal adder_s_net_x4: std_logic_vector(19 downto 0);
  signal adder_s_net_x5: std_logic_vector(19 downto 0);
  signal adder_s_net_x6: std_logic_vector(19 downto 0);
  signal adder_s_net_x7: std_logic_vector(19 downto 0);
  signal ce_1_sg_x76: std_logic;
  signal clk_1_sg_x76: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  ce_1_sg_x76 <= ce_1;
  clk_1_sg_x76 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_e395239523: entity work.bussify_entity_c32f93b775
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_254c41df9c: entity work.conv1_entity_254c41df9c
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_170b394fa6: entity work.conv1_entity_254c41df9c
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_ffbee01946: entity work.conv1_entity_254c41df9c
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_8d4be2e173: entity work.conv1_entity_254c41df9c
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_edfe8ef4dd: entity work.debus_entity_9e67f505ae
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_relational/a_debus"

entity a_debus_entity_019babc48f is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    msb_lsb_out1: out std_logic_vector(3 downto 0)
  );
end a_debus_entity_019babc48f;

architecture structural of a_debus_entity_019babc48f is
  signal constant_op_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net: std_logic_vector(3 downto 0);

begin
  constant_op_net_x0 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x0;

  reinterpret1: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 4,
      y_width => 4
    )
    port map (
      x => constant_op_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_relational"

entity bus_relational_entity_ea2675d756 is
  port (
    a: in std_logic_vector(3 downto 0); 
    b: in std_logic_vector(3 downto 0); 
    a_b: out std_logic
  );
end bus_relational_entity_ea2675d756;

architecture structural of bus_relational_entity_ea2675d756 is
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic;
  signal reinterpret_out_output_port_net_x1: std_logic_vector(3 downto 0);
  signal relational1_op_net_x0: std_logic;

begin
  constant_op_net_x1 <= a;
  reinterpret_out_output_port_net_x1 <= b;
  a_b <= reinterpret1_output_port_net_x3;

  a_debus_019babc48f: entity work.a_debus_entity_019babc48f
    port map (
      bus_in => constant_op_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  b_debus_7952c3e710: entity work.a_debus_entity_019babc48f
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  bussify_df4eac8774: entity work.bussify_entity_ad099992fc
    port map (
      in1 => relational1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x3
    );

  relational1: entity work.relational_d930162434
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/bus_sub"

entity bus_sub_entity_2680215111 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(37 downto 0)
  );
end bus_sub_entity_2680215111;

architecture structural of bus_sub_entity_2680215111 is
  signal addsub1_s_net_x0: std_logic_vector(18 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(18 downto 0);
  signal ce_1_sg_x77: std_logic;
  signal clk_1_sg_x77: std_logic;
  signal concatenate_y_net_x4: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(37 downto 0);
  signal dmux0_q_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x4 <= a;
  dmux0_q_net_x3 <= b;
  ce_1_sg_x77 <= ce_1;
  clk_1_sg_x77 <= clk_1;
  dout <= concatenate_y_net_x5;

  a_debus_af86cbcf92: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_c9b173d075a3b6d7",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 18,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 19,
      core_name0 => "addsb_11_0_c9b173d075a3b6d7",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 19,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_b879dc1045: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => dmux0_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_8231241e68: entity work.op_bussify_entity_a6d4bedd3c
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/munge/join"

entity join_entity_3e6265795f is
  port (
    in1: in std_logic_vector(1 downto 0); 
    in2: in std_logic_vector(1 downto 0); 
    bus_out: out std_logic_vector(3 downto 0)
  );
end join_entity_3e6265795f;

architecture structural of join_entity_3e6265795f is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(1 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(1 downto 0);

begin
  reinterpret2_output_port_net_x1 <= in1;
  reinterpret1_output_port_net_x1 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x1,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret1_output_port_net_x1,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/munge/split"

entity split_entity_eadf33f9d0 is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    lsb_out1: out std_logic_vector(1 downto 0); 
    msb_out2: out std_logic_vector(1 downto 0)
  );
end split_entity_eadf33f9d0;

architecture structural of split_entity_eadf33f9d0 is
  signal reinterpret1_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net: std_logic_vector(1 downto 0);
  signal slice2_y_net: std_logic_vector(1 downto 0);

begin
  reinterpret_output_port_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out2 <= reinterpret2_output_port_net_x2;

  reinterpret1: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_9a54e08c7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => reinterpret_output_port_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => reinterpret_output_port_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/munge"

entity munge_entity_8c0725027d is
  port (
    din: in std_logic_vector(3 downto 0); 
    dout: out std_logic_vector(3 downto 0)
  );
end munge_entity_8c0725027d;

architecture structural of munge_entity_8c0725027d is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(3 downto 0);

begin
  concatenate_y_net_x6 <= din;
  dout <= reinterpret_out_output_port_net_x2;

  join_3e6265795f: entity work.join_entity_3e6265795f
    port map (
      in1 => reinterpret2_output_port_net_x2,
      in2 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x0
    );

  reinterpret: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x6,
      output_port => reinterpret_output_port_net_x0
    );

  reinterpret_out: entity work.reinterpret_d610556e85
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concatenate_y_net_x0,
      output_port => reinterpret_out_output_port_net_x2
    );

  split_eadf33f9d0: entity work.split_entity_eadf33f9d0
    port map (
      bus_in => reinterpret_output_port_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/mux/d_bussify"

entity d_bussify_entity_815212a6f1 is
  port (
    in1: in std_logic_vector(19 downto 0); 
    in2: in std_logic_vector(19 downto 0); 
    in3: in std_logic_vector(19 downto 0); 
    in4: in std_logic_vector(19 downto 0); 
    bus_out: out std_logic_vector(79 downto 0)
  );
end d_bussify_entity_815212a6f1;

architecture structural of d_bussify_entity_815212a6f1 is
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal mux0_y_net_x0: std_logic_vector(19 downto 0);
  signal mux1_y_net_x0: std_logic_vector(19 downto 0);
  signal mux2_y_net_x0: std_logic_vector(19 downto 0);
  signal mux3_y_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(19 downto 0);

begin
  mux0_y_net_x0 <= in1;
  mux1_y_net_x0 <= in2;
  mux2_y_net_x0 <= in3;
  mux3_y_net_x0 <= in4;
  bus_out <= concatenate_y_net_x4;

  concatenate: entity work.concat_f86ebb6084
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x4
    );

  reinterpret1: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux0_y_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux1_y_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux2_y_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux3_y_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/mux/expand0"

entity expand0_entity_2b461ef222 is
  port (
    bus_in: in std_logic_vector(79 downto 0); 
    lsb_out1: out std_logic_vector(19 downto 0); 
    msb_out4: out std_logic_vector(19 downto 0); 
    out2: out std_logic_vector(19 downto 0); 
    out3: out std_logic_vector(19 downto 0)
  );
end expand0_entity_2b461ef222;

architecture structural of expand0_entity_2b461ef222 is
  signal concatenate_y_net_x2: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic_vector(19 downto 0);
  signal slice2_y_net: std_logic_vector(19 downto 0);
  signal slice3_y_net: std_logic_vector(19 downto 0);
  signal slice4_y_net: std_logic_vector(19 downto 0);

begin
  concatenate_y_net_x2 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_713b6c5d29
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 19,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 39,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 59,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 79,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/mux/sel_expand"

entity sel_expand_entity_41b2560930 is
  port (
    bus_in: in std_logic_vector(3 downto 0); 
    lsb_out1: out std_logic; 
    msb_out4: out std_logic; 
    out2: out std_logic; 
    out3: out std_logic
  );
end sel_expand_entity_41b2560930;

architecture structural of sel_expand_entity_41b2560930 is
  signal concatenate_y_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic;
  signal reinterpret3_output_port_net_x0: std_logic;
  signal reinterpret4_output_port_net_x0: std_logic;
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic;
  signal slice3_y_net: std_logic;
  signal slice4_y_net: std_logic;

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_81130c7f2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => slice1_y_net,
      output_port(0) => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_81130c7f2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => slice2_y_net,
      output_port(0) => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_81130c7f2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => slice3_y_net,
      output_port(0) => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_81130c7f2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => slice4_y_net,
      output_port(0) => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/mux"

entity mux_entity_e2fd897480 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d0: in std_logic_vector(79 downto 0); 
    d1: in std_logic_vector(79 downto 0); 
    sel: in std_logic_vector(3 downto 0); 
    out_x0: out std_logic_vector(79 downto 0)
  );
end mux_entity_e2fd897480;

architecture structural of mux_entity_e2fd897480 is
  signal ce_1_sg_x78: std_logic;
  signal clk_1_sg_x78: std_logic;
  signal concatenate_y_net_x6: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(79 downto 0);
  signal mux0_y_net_x0: std_logic_vector(19 downto 0);
  signal mux1_y_net_x0: std_logic_vector(19 downto 0);
  signal mux2_y_net_x0: std_logic_vector(19 downto 0);
  signal mux3_y_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic;
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic;
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic;

begin
  ce_1_sg_x78 <= ce_1;
  clk_1_sg_x78 <= clk_1;
  concatenate_y_net_x6 <= d0;
  concatenate_y_net_x7 <= d1;
  concatenate_y_net_x8 <= sel;
  out_x0 <= concatenate_y_net_x9;

  d_bussify_815212a6f1: entity work.d_bussify_entity_815212a6f1
    port map (
      in1 => mux0_y_net_x0,
      in2 => mux1_y_net_x0,
      in3 => mux2_y_net_x0,
      in4 => mux3_y_net_x0,
      bus_out => concatenate_y_net_x9
    );

  expand0_2b461ef222: entity work.expand0_entity_2b461ef222
    port map (
      bus_in => concatenate_y_net_x6,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  expand1_559314c247: entity work.expand0_entity_2b461ef222
    port map (
      bus_in => concatenate_y_net_x7,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

  mux0: entity work.mux_ce20fdf7b8
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      d0 => reinterpret4_output_port_net_x0,
      d1 => reinterpret4_output_port_net_x1,
      sel(0) => reinterpret4_output_port_net_x2,
      y => mux0_y_net_x0
    );

  mux1: entity work.mux_ce20fdf7b8
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      d0 => reinterpret3_output_port_net_x0,
      d1 => reinterpret3_output_port_net_x1,
      sel(0) => reinterpret3_output_port_net_x2,
      y => mux1_y_net_x0
    );

  mux2: entity work.mux_ce20fdf7b8
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      d0 => reinterpret2_output_port_net_x0,
      d1 => reinterpret2_output_port_net_x1,
      sel(0) => reinterpret2_output_port_net_x2,
      y => mux2_y_net_x0
    );

  mux3: entity work.mux_ce20fdf7b8
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      d0 => reinterpret1_output_port_net_x0,
      d1 => reinterpret1_output_port_net_x1,
      sel(0) => reinterpret1_output_port_net_x2,
      y => mux3_y_net_x0
    );

  sel_expand_41b2560930: entity work.sel_expand_entity_41b2560930
    port map (
      bus_in => concatenate_y_net_x8,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct/shift_replicate"

entity shift_replicate_entity_a296056610 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic_vector(3 downto 0)
  );
end shift_replicate_entity_a296056610;

architecture structural of shift_replicate_entity_a296056610 is
  signal ce_1_sg_x79: std_logic;
  signal clk_1_sg_x79: std_logic;
  signal concatenate_y_net_x10: std_logic_vector(3 downto 0);
  signal din0_0_q_net_x0: std_logic;
  signal din0_1_q_net_x0: std_logic;
  signal din0_2_q_net_x0: std_logic;
  signal din0_3_q_net_x0: std_logic;
  signal slice0_y_net_x0: std_logic;

begin
  ce_1_sg_x79 <= ce_1;
  clk_1_sg_x79 <= clk_1;
  slice0_y_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x10;

  bussify_3fc834941b: entity work.bussify_entity_6bd38bcd1d
    port map (
      in1 => din0_0_q_net_x0,
      in2 => din0_1_q_net_x0,
      in3 => din0_2_q_net_x0,
      in4 => din0_3_q_net_x0,
      bus_out => concatenate_y_net_x10
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => slice0_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_0_q_net_x0
    );

  din0_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => slice0_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_1_q_net_x0
    );

  din0_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => slice0_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_2_q_net_x0
    );

  din0_3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x79,
      clk => clk_1_sg_x79,
      d(0) => slice0_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => din0_3_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/butterfly_direct"

entity butterfly_direct_entity_63ba888001 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_63ba888001;

architecture structural of butterfly_direct_entity_63ba888001 is
  signal ce_1_sg_x80: std_logic;
  signal clk_1_sg_x80: std_logic;
  signal concat_y_net_x3: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x13: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x4: std_logic_vector(35 downto 0);
  signal mux_y_net_x0: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;

begin
  concatenate_y_net_x13 <= a;
  dmux0_q_net_x4 <= b;
  ce_1_sg_x80 <= ce_1;
  clk_1_sg_x80 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x0 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x5;
  sync_out <= delay0_q_net_x0;

  bus_add_a60c7dc670: entity work.bus_add_entity_a60c7dc670
    port map (
      a => concatenate_y_net_x13,
      b => dmux0_q_net_x4,
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      dout => concatenate_y_net_x3
    );

  bus_convert_7b742cca79: entity work.bus_convert_entity_7b742cca79
    port map (
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_f69635d38b: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_74bb60a7d0: entity work.bus_norm0_entity_74bb60a7d0
    port map (
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_b00e4bc012: entity work.bus_norm1_entity_b00e4bc012
    port map (
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_ea2675d756: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x5
    );

  bus_scale_af5b203396: entity work.bus_scale_entity_316a2a993e
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_2680215111: entity work.bus_sub_entity_2680215111
    port map (
      a => concatenate_y_net_x13,
      b => dmux0_q_net_x4,
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_4822199898
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x80,
      clk => clk_1_sg_x80,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => delay0_q_net_x0
    );

  munge_8c0725027d: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_e2fd897480: entity work.mux_entity_e2fd897480
    port map (
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_a296056610: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x80,
      clk_1 => clk_1_sg_x80,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/debus_addr"

entity debus_addr_entity_47d8ecebba is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(11 downto 0); 
    msb_out3: out std_logic_vector(11 downto 0); 
    out2: out std_logic_vector(11 downto 0)
  );
end debus_addr_entity_47d8ecebba;

architecture structural of debus_addr_entity_47d8ecebba is
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(11 downto 0);
  signal slice1_y_net: std_logic_vector(11 downto 0);
  signal slice2_y_net: std_logic_vector(11 downto 0);
  signal slice3_y_net: std_logic_vector(11 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out3 <= reinterpret3_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 36,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 23,
      x_width => 36,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 35,
      x_width => 36,
      y_width => 12
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/debus_we"

entity debus_we_entity_ddd27e7170 is
  port (
    bus_in: in std_logic_vector(2 downto 0); 
    lsb_out1: out std_logic; 
    msb_out3: out std_logic; 
    out2: out std_logic
  );
end debus_we_entity_ddd27e7170;

architecture structural of debus_we_entity_ddd27e7170 is
  signal concatenate_y_net_x0: std_logic_vector(2 downto 0);
  signal slice1_y_net_x0: std_logic;
  signal slice2_y_net_x0: std_logic;
  signal slice3_y_net_x0: std_logic;

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= slice1_y_net_x0;
  msb_out3 <= slice3_y_net_x0;
  out2 <= slice2_y_net_x0;

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice1_y_net_x0
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice2_y_net_x0
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => concatenate_y_net_x0,
      y(0) => slice3_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/rep_addr/bussify"

entity bussify_entity_1f1b293ba3 is
  port (
    in1: in std_logic_vector(11 downto 0); 
    in2: in std_logic_vector(11 downto 0); 
    in3: in std_logic_vector(11 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end bussify_entity_1f1b293ba3;

architecture structural of bussify_entity_1f1b293ba3 is
  signal concatenate_y_net_x1: std_logic_vector(35 downto 0);
  signal din3_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_2_q_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(11 downto 0);

begin
  din3_0_q_net_x0 <= in1;
  din3_1_q_net_x0 <= in2;
  din3_2_q_net_x0 <= in3;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_d7d801964d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_0_q_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_1_q_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_75275f6c4a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din3_2_q_net_x0,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/rep_addr"

entity rep_addr_entity_b150ee5367 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(35 downto 0)
  );
end rep_addr_entity_b150ee5367;

architecture structural of rep_addr_entity_b150ee5367 is
  signal addr0_op_net_x0: std_logic_vector(11 downto 0);
  signal ce_1_sg_x81: std_logic;
  signal clk_1_sg_x81: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal din0_0_q_net: std_logic_vector(11 downto 0);
  signal din1_0_q_net: std_logic_vector(11 downto 0);
  signal din1_1_q_net: std_logic_vector(11 downto 0);
  signal din2_0_q_net: std_logic_vector(11 downto 0);
  signal din2_1_q_net: std_logic_vector(11 downto 0);
  signal din2_2_q_net: std_logic_vector(11 downto 0);
  signal din3_0_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_1_q_net_x0: std_logic_vector(11 downto 0);
  signal din3_2_q_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x81 <= ce_1;
  clk_1_sg_x81 <= clk_1;
  addr0_op_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_1f1b293ba3: entity work.bussify_entity_1f1b293ba3
    port map (
      in1 => din3_0_q_net_x0,
      in2 => din3_1_q_net_x0,
      in3 => din3_2_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => addr0_op_net_x0,
      en => '1',
      rst => '1',
      q => din0_0_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_0_q_net
    );

  din1_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_1_q_net
    );

  din2_0: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      clr => '0',
      d => din1_0_q_net,
      q => din2_0_q_net
    );

  din2_1: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      clr => '0',
      d => din1_1_q_net,
      q => din2_1_q_net
    );

  din2_2: entity work.delay_87cc993d41
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      clr => '0',
      d => din1_0_q_net,
      q => din2_2_q_net
    );

  din3_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => din2_0_q_net,
      en => '1',
      rst => '1',
      q => din3_0_q_net_x0
    );

  din3_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => din2_1_q_net,
      en => '1',
      rst => '1',
      q => din3_1_q_net_x0
    );

  din3_2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      d => din2_2_q_net,
      en => '1',
      rst => '1',
      q => din3_2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/rep_we/bussify"

entity bussify_entity_f6b3da5312 is
  port (
    in1: in std_logic; 
    in2: in std_logic; 
    in3: in std_logic; 
    bus_out: out std_logic_vector(2 downto 0)
  );
end bussify_entity_f6b3da5312;

architecture structural of bussify_entity_f6b3da5312 is
  signal concatenate_y_net_x1: std_logic_vector(2 downto 0);
  signal din3_0_q_net_x0: std_logic;
  signal din3_1_q_net_x0: std_logic;
  signal din3_2_q_net_x0: std_logic;
  signal reinterpret1_output_port_net: std_logic;
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic;

begin
  din3_0_q_net_x0 <= in1;
  din3_1_q_net_x0 <= in2;
  din3_2_q_net_x0 <= in3;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_452c4d3410
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2(0) => reinterpret3_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_0_q_net_x0,
      output_port(0) => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_1_q_net_x0,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => din3_2_q_net_x0,
      output_port(0) => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0/rep_we"

entity rep_we_entity_41df2e67d6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic_vector(2 downto 0)
  );
end rep_we_entity_41df2e67d6;

architecture structural of rep_we_entity_41df2e67d6 is
  signal ce_1_sg_x82: std_logic;
  signal clk_1_sg_x82: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(2 downto 0);
  signal din0_0_q_net: std_logic;
  signal din1_0_q_net: std_logic;
  signal din1_1_q_net: std_logic;
  signal din2_0_q_net: std_logic;
  signal din2_1_q_net: std_logic;
  signal din2_2_q_net: std_logic;
  signal din3_0_q_net_x0: std_logic;
  signal din3_1_q_net_x0: std_logic;
  signal din3_2_q_net_x0: std_logic;
  signal we0_op_net_x0: std_logic;

begin
  ce_1_sg_x82 <= ce_1;
  clk_1_sg_x82 <= clk_1;
  we0_op_net_x0 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_f6b3da5312: entity work.bussify_entity_f6b3da5312
    port map (
      in1 => din3_0_q_net_x0,
      in2 => din3_1_q_net_x0,
      in3 => din3_2_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => we0_op_net_x0,
      q(0) => din0_0_q_net
    );

  din1_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din0_0_q_net,
      q(0) => din1_0_q_net
    );

  din1_1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din0_0_q_net,
      q(0) => din1_1_q_net
    );

  din2_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din1_0_q_net,
      q(0) => din2_0_q_net
    );

  din2_1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din1_1_q_net,
      q(0) => din2_1_q_net
    );

  din2_2: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din1_0_q_net,
      q(0) => din2_2_q_net
    );

  din3_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din2_0_q_net,
      q(0) => din3_0_q_net_x0
    );

  din3_1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din2_1_q_net,
      q(0) => din3_1_q_net_x0
    );

  din3_2: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x82,
      clk => clk_1_sg_x82,
      clr => '0',
      d(0) => din2_2_q_net,
      q(0) => din3_2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1/delay0"

entity delay0_entity_bcdc7ba653 is
  port (
    addr: in std_logic_vector(11 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    we: in std_logic; 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_bcdc7ba653;

architecture structural of delay0_entity_bcdc7ba653 is
  signal addr0_op_net_x1: std_logic_vector(11 downto 0);
  signal bram0_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram4_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram5_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram6_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram7_data_out_net_x0: std_logic_vector(3 downto 0);
  signal bram8_data_out_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x83: std_logic;
  signal clk_1_sg_x83: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(2 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(35 downto 0);
  signal ddin_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(3 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret5_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret6_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret7_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret8_output_port_net_x0: std_logic_vector(3 downto 0);
  signal reinterpret9_output_port_net_x0: std_logic_vector(3 downto 0);
  signal slice1_y_net_x0: std_logic;
  signal slice2_y_net_x0: std_logic;
  signal slice3_y_net_x0: std_logic;
  signal we0_op_net_x1: std_logic;

begin
  addr0_op_net_x1 <= addr;
  ce_1_sg_x83 <= ce_1;
  clk_1_sg_x83 <= clk_1;
  reinterpret1_output_port_net_x2 <= din;
  we0_op_net_x1 <= we;
  dout <= concatenate_y_net_x4;

  bram0: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret3_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret9_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice3_y_net_x0,
      data_out => bram0_data_out_net_x0
    );

  bram1: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret2_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret8_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice2_y_net_x0,
      data_out => bram1_data_out_net_x0
    );

  bram2: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret7_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram2_data_out_net_x0
    );

  bram3: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret3_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret6_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice3_y_net_x0,
      data_out => bram3_data_out_net_x0
    );

  bram4: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret2_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret5_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice2_y_net_x0,
      data_out => bram4_data_out_net_x0
    );

  bram5: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret4_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram5_data_out_net_x0
    );

  bram6: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret3_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret3_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice3_y_net_x0,
      data_out => bram6_data_out_net_x0
    );

  bram7: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret2_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret2_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice2_y_net_x0,
      data_out => bram7_data_out_net_x0
    );

  bram8: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 12,
      c_width => 4,
      core_name0 => "bmg_72_fa6496d84f038019",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      data_in => reinterpret1_output_port_net_x1,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram8_data_out_net_x0
    );

  ddin: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x83,
      clk => clk_1_sg_x83,
      clr => '0',
      d => reinterpret1_output_port_net_x2,
      q => ddin_q_net_x0
    );

  debus_addr_47d8ecebba: entity work.debus_addr_entity_47d8ecebba
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out3 => reinterpret3_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0
    );

  debus_din_cf53163a90: entity work.debus_din_entity_d2fe8dc95c
    port map (
      bus_in => ddin_q_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out9 => reinterpret9_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1,
      out4 => reinterpret4_output_port_net_x0,
      out5 => reinterpret5_output_port_net_x0,
      out6 => reinterpret6_output_port_net_x0,
      out7 => reinterpret7_output_port_net_x0,
      out8 => reinterpret8_output_port_net_x0
    );

  debus_we_ddd27e7170: entity work.debus_we_entity_ddd27e7170
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => slice1_y_net_x0,
      msb_out3 => slice3_y_net_x0,
      out2 => slice2_y_net_x0
    );

  din_bussify_59bda723ef: entity work.din_bussify_entity_e936a8b4d0
    port map (
      in1 => bram0_data_out_net_x0,
      in2 => bram1_data_out_net_x0,
      in3 => bram2_data_out_net_x0,
      in4 => bram3_data_out_net_x0,
      in5 => bram4_data_out_net_x0,
      in6 => bram5_data_out_net_x0,
      in7 => bram6_data_out_net_x0,
      in8 => bram7_data_out_net_x0,
      in9 => bram8_data_out_net_x0,
      bus_out => concatenate_y_net_x4
    );

  rep_addr_b150ee5367: entity work.rep_addr_entity_b150ee5367
    port map (
      ce_1 => ce_1_sg_x83,
      clk_1 => clk_1_sg_x83,
      in_x0 => addr0_op_net_x1,
      out_x0 => concatenate_y_net_x2
    );

  rep_we_41df2e67d6: entity work.rep_we_entity_41df2e67d6
    port map (
      ce_1 => ce_1_sg_x83,
      clk_1 => clk_1_sg_x83,
      in_x0 => we0_op_net_x1,
      out_x0 => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_1"

entity fft_stage_1_entity_f280a22ded is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_1_entity_f280a22ded;

architecture structural of fft_stage_1_entity_f280a22ded is
  signal addr0_op_net_x1: std_logic_vector(11 downto 0);
  signal addr1_op_net_x1: std_logic_vector(11 downto 0);
  signal ce_1_sg_x88: std_logic;
  signal clk_1_sg_x88: std_logic;
  signal concatenate_y_net_x15: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(35 downto 0);
  signal constant_op_net_x0: std_logic;
  signal counter_op_net: std_logic_vector(12 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din1_q_net: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x4: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal dsync2_q_net: std_logic;
  signal fft_shift_net_x0: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;
  signal sync_net_x0: std_logic;
  signal we0_op_net_x1: std_logic;
  signal we1_op_net_x1: std_logic;

begin
  ce_1_sg_x88 <= ce_1;
  clk_1_sg_x88 <= clk_1;
  reinterpret1_output_port_net_x0 <= in1;
  reinterpret1_output_port_net_x6 <= in2;
  constant_op_net_x0 <= of_in;
  fft_shift_net_x0 <= shift;
  sync_net_x0 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x7;
  sync_out <= delay0_q_net_x1;

  addr0: entity work.counter_6cd08a247e
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      op => addr0_op_net_x1
    );

  addr1: entity work.counter_6cd08a247e
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      op => addr1_op_net_x1
    );

  butterfly_direct_63ba888001: entity work.butterfly_direct_entity_63ba888001
    port map (
      a => concatenate_y_net_x15,
      b => dmux0_q_net_x4,
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x1,
      a_bw => reinterpret1_output_port_net_x7,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x5,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.counter_c48d6dcab5
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      rst(0) => dsync2_q_net,
      op => counter_op_net
    );

  delay0_bcdc7ba653: entity work.delay0_entity_bcdc7ba653
    port map (
      addr => addr0_op_net_x1,
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      din => reinterpret1_output_port_net_x6,
      we => we0_op_net_x1,
      dout => concatenate_y_net_x4
    );

  delay1_d0e0aa0b30: entity work.delay0_entity_bcdc7ba653
    port map (
      addr => addr1_op_net_x1,
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      din => mux1_y_net_x0,
      we => we1_op_net_x1,
      dout => concatenate_y_net_x15
    );

  din0: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => din0_q_net
    );

  din1: entity work.delay_4b00a70dea
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d => din0_q_net,
      q => din1_q_net
    );

  dmux0: entity work.delay_1b04a69dde
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x4
    );

  dsync0: entity work.delay_c53de546ea
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d(0) => sync_net_x0,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_14a6a51cbc
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d(0) => dsync2_q_net,
      q(0) => dsync1_q_net_x0
    );

  dsync2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync2_q_net
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x5,
      d1(0) => constant_op_net_x0,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d0 => concatenate_y_net_x4,
      d1 => din1_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x88,
      clk => clk_1_sg_x88,
      clr => '0',
      d0 => din1_q_net,
      d1 => concatenate_y_net_x4,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x0,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 13,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_c758427ca8: entity work.sync_delay_entity_c43fa8c0d9
    port map (
      ce_1 => ce_1_sg_x88,
      clk_1 => clk_1_sg_x88,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x1
    );

  we0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => we0_op_net_x1
    );

  we1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => we1_op_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_add/b_debus"

entity b_debus_entity_97187af928 is
  port (
    bus_in: in std_logic_vector(37 downto 0); 
    lsb_out1: out std_logic_vector(18 downto 0); 
    msb_out2: out std_logic_vector(18 downto 0)
  );
end b_debus_entity_97187af928;

architecture structural of b_debus_entity_97187af928 is
  signal concatenate_y_net_x0: std_logic_vector(37 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(18 downto 0);
  signal slice1_y_net: std_logic_vector(18 downto 0);
  signal slice2_y_net: std_logic_vector(18 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_63700884f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 18,
      x_width => 38,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 37,
      x_width => 38,
      y_width => 19
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_add/op_bussify"

entity op_bussify_entity_cf1986e0b4 is
  port (
    in1: in std_logic_vector(19 downto 0); 
    in2: in std_logic_vector(19 downto 0); 
    bus_out: out std_logic_vector(39 downto 0)
  );
end op_bussify_entity_cf1986e0b4;

architecture structural of op_bussify_entity_cf1986e0b4 is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(19 downto 0);

begin
  addsub1_s_net_x0 <= in1;
  addsub2_s_net_x0 <= in2;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_9e724c4b50
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub1_s_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => addsub2_s_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_add"

entity bus_add_entity_277738c818 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(37 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(39 downto 0)
  );
end bus_add_entity_277738c818;

architecture structural of bus_add_entity_277738c818 is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal ce_1_sg_x89: std_logic;
  signal clk_1_sg_x89: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  reinterpret1_output_port_net_x3 <= a;
  concatenate_y_net_x2 <= b;
  ce_1_sg_x89 <= ce_1;
  clk_1_sg_x89 <= clk_1;
  dout <= concatenate_y_net_x3;

  a_debus_08d3df532c: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_6bbb8fb0d8f20abe",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x89,
      clk => clk_1_sg_x89,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_6bbb8fb0d8f20abe",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret1_output_port_net_x2,
      b => reinterpret1_output_port_net_x0,
      ce => ce_1_sg_x89,
      clk => clk_1_sg_x89,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_97187af928: entity work.b_debus_entity_97187af928
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_cf1986e0b4: entity work.op_bussify_entity_cf1986e0b4
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_convert/conv1/convert"

entity convert_entity_8b4a784542 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(20 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end convert_entity_8b4a784542;

architecture structural of convert_entity_8b4a784542 is
  signal adder_s_net_x4: std_logic_vector(17 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x90: std_logic;
  signal clk_1_sg_x90: std_logic;
  signal concat_y_net: std_logic_vector(21 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(21 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(20 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x90 <= ce_1;
  clk_1_sg_x90 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 19,
      a_width => 22,
      b_arith => xlUnsigned,
      b_bin_pt => 19,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 23,
      core_name0 => "addsb_11_0_1f22b9fac024cf00",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 23,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 18
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      clr => '0',
      en => "1",
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_4709ea49b5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_e6bc20c81b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_c84451c80b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_convert/conv1"

entity conv1_entity_f8f57d1952 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(20 downto 0); 
    dout: out std_logic_vector(17 downto 0); 
    of_x0: out std_logic
  );
end conv1_entity_f8f57d1952;

architecture structural of conv1_entity_f8f57d1952 is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal all_0s_y_net: std_logic;
  signal all_1s_y_net: std_logic;
  signal and_y_net_x0: std_logic;
  signal ce_1_sg_x91: std_logic;
  signal clk_1_sg_x91: std_logic;
  signal invert1_op_net: std_logic;
  signal invert2_op_net: std_logic;
  signal invert3_op_net: std_logic;
  signal reinterpret4_output_port_net_x1: std_logic_vector(20 downto 0);
  signal slice1_y_net: std_logic;
  signal slice2_y_net: std_logic;
  signal slice3_y_net: std_logic;

begin
  ce_1_sg_x91 <= ce_1;
  clk_1_sg_x91 <= clk_1;
  reinterpret4_output_port_net_x1 <= din;
  dout <= adder_s_net_x5;
  of_x0 <= and_y_net_x0;

  all_0s: entity work.logical_fe87bb6ae4
    port map (
      ce => ce_1_sg_x91,
      clk => clk_1_sg_x91,
      clr => '0',
      d0(0) => invert1_op_net,
      d1(0) => invert2_op_net,
      d2(0) => invert3_op_net,
      y(0) => all_0s_y_net
    );

  all_1s: entity work.logical_fe87bb6ae4
    port map (
      ce => ce_1_sg_x91,
      clk => clk_1_sg_x91,
      clr => '0',
      d0(0) => slice1_y_net,
      d1(0) => slice2_y_net,
      d2(0) => slice3_y_net,
      y(0) => all_1s_y_net
    );

  and_x0: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => all_0s_y_net,
      d1(0) => all_1s_y_net,
      y(0) => and_y_net_x0
    );

  convert_8b4a784542: entity work.convert_entity_8b4a784542
    port map (
      ce_1 => ce_1_sg_x91,
      clk_1 => clk_1_sg_x91,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  invert1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x91,
      clk => clk_1_sg_x91,
      clr => '0',
      ip(0) => slice1_y_net,
      op(0) => invert1_op_net
    );

  invert2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x91,
      clk => clk_1_sg_x91,
      clr => '0',
      ip(0) => slice2_y_net,
      op(0) => invert2_op_net
    );

  invert3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x91,
      clk => clk_1_sg_x91,
      clr => '0',
      ip(0) => slice3_y_net,
      op(0) => invert3_op_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 20,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 19,
      new_msb => 19,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 18,
      x_width => 21,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x1,
      y(0) => slice3_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_convert/debus"

entity debus_entity_0c420b862c is
  port (
    bus_in: in std_logic_vector(83 downto 0); 
    lsb_out1: out std_logic_vector(20 downto 0); 
    msb_out4: out std_logic_vector(20 downto 0); 
    out2: out std_logic_vector(20 downto 0); 
    out3: out std_logic_vector(20 downto 0)
  );
end debus_entity_0c420b862c;

architecture structural of debus_entity_0c420b862c is
  signal concatenate_y_net_x0: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(20 downto 0);
  signal slice1_y_net: std_logic_vector(20 downto 0);
  signal slice2_y_net: std_logic_vector(20 downto 0);
  signal slice3_y_net: std_logic_vector(20 downto 0);
  signal slice4_y_net: std_logic_vector(20 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out4 <= reinterpret4_output_port_net_x2;
  out2 <= reinterpret2_output_port_net_x2;
  out3 <= reinterpret3_output_port_net_x2;

  reinterpret1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  reinterpret3: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x2
    );

  reinterpret4: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 20,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 21,
      new_msb => 41,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 42,
      new_msb => 62,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 63,
      new_msb => 83,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_convert"

entity bus_convert_entity_43c000ec6d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(83 downto 0); 
    dout: out std_logic_vector(71 downto 0); 
    overflow: out std_logic_vector(3 downto 0)
  );
end bus_convert_entity_43c000ec6d;

architecture structural of bus_convert_entity_43c000ec6d is
  signal adder_s_net_x5: std_logic_vector(17 downto 0);
  signal adder_s_net_x6: std_logic_vector(17 downto 0);
  signal adder_s_net_x7: std_logic_vector(17 downto 0);
  signal adder_s_net_x8: std_logic_vector(17 downto 0);
  signal and_y_net_x4: std_logic;
  signal and_y_net_x5: std_logic;
  signal and_y_net_x6: std_logic;
  signal and_y_net_x7: std_logic;
  signal ce_1_sg_x98: std_logic;
  signal clk_1_sg_x98: std_logic;
  signal concatenate_y_net_x3: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(3 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic_vector(20 downto 0);

begin
  ce_1_sg_x98 <= ce_1;
  clk_1_sg_x98 <= clk_1;
  concatenate_y_net_x3 <= din;
  dout <= concatenate_y_net_x4;
  overflow <= concatenate_y_net_x5;

  bussify_19c1e8b1e1: entity work.bussify_entity_904656ce6f
    port map (
      in1 => adder_s_net_x5,
      in2 => adder_s_net_x6,
      in3 => adder_s_net_x7,
      in4 => adder_s_net_x8,
      bus_out => concatenate_y_net_x4
    );

  conv1_f8f57d1952: entity work.conv1_entity_f8f57d1952
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      din => reinterpret4_output_port_net_x2,
      dout => adder_s_net_x5,
      of_x0 => and_y_net_x4
    );

  conv2_cd18bf91b1: entity work.conv1_entity_f8f57d1952
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      din => reinterpret3_output_port_net_x2,
      dout => adder_s_net_x6,
      of_x0 => and_y_net_x5
    );

  conv3_a19e34497a: entity work.conv1_entity_f8f57d1952
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      din => reinterpret2_output_port_net_x2,
      dout => adder_s_net_x7,
      of_x0 => and_y_net_x6
    );

  conv4_eba6811c4d: entity work.conv1_entity_f8f57d1952
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      din => reinterpret1_output_port_net_x2,
      dout => adder_s_net_x8,
      of_x0 => and_y_net_x7
    );

  debus_0c420b862c: entity work.debus_entity_0c420b862c
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

  of_bussify_691c7fc8cf: entity work.bussify_entity_6bd38bcd1d
    port map (
      in1 => and_y_net_x4,
      in2 => and_y_net_x5,
      in3 => and_y_net_x6,
      in4 => and_y_net_x7,
      bus_out => concatenate_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_norm0/bussify"

entity bussify_entity_83bee71966 is
  port (
    in1: in std_logic_vector(20 downto 0); 
    in2: in std_logic_vector(20 downto 0); 
    in3: in std_logic_vector(20 downto 0); 
    in4: in std_logic_vector(20 downto 0); 
    bus_out: out std_logic_vector(83 downto 0)
  );
end bussify_entity_83bee71966;

architecture structural of bussify_entity_83bee71966 is
  signal concatenate_y_net_x0: std_logic_vector(83 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(20 downto 0);

begin
  conv1_dout_net_x0 <= in1;
  conv2_dout_net_x0 <= in2;
  conv3_dout_net_x0 <= in3;
  conv4_dout_net_x0 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_356a264444
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv1_dout_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv2_dout_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv3_dout_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_f0ca8483cb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => conv4_dout_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_norm0/debus"

entity debus_entity_fe21c1b916 is
  port (
    bus_in: in std_logic_vector(79 downto 0); 
    lsb_out1: out std_logic_vector(19 downto 0); 
    msb_out4: out std_logic_vector(19 downto 0); 
    out2: out std_logic_vector(19 downto 0); 
    out3: out std_logic_vector(19 downto 0)
  );
end debus_entity_fe21c1b916;

architecture structural of debus_entity_fe21c1b916 is
  signal concat_y_net_x0: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal slice1_y_net: std_logic_vector(19 downto 0);
  signal slice2_y_net: std_logic_vector(19 downto 0);
  signal slice3_y_net: std_logic_vector(19 downto 0);
  signal slice4_y_net: std_logic_vector(19 downto 0);

begin
  concat_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_f661f8d9b7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 19,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 20,
      new_msb => 39,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 59,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 60,
      new_msb => 79,
      x_width => 80,
      y_width => 20
    )
    port map (
      x => concat_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_norm0"

entity bus_norm0_entity_376e099b6a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(83 downto 0)
  );
end bus_norm0_entity_376e099b6a;

architecture structural of bus_norm0_entity_376e099b6a is
  signal ce_1_sg_x99: std_logic;
  signal clk_1_sg_x99: std_logic;
  signal concat_y_net_x1: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(83 downto 0);
  signal conv1_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv2_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv3_dout_net_x0: std_logic_vector(20 downto 0);
  signal conv4_dout_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x99 <= ce_1;
  clk_1_sg_x99 <= clk_1;
  concat_y_net_x1 <= din;
  dout <= concatenate_y_net_x1;

  bussify_83bee71966: entity work.bussify_entity_83bee71966
    port map (
      in1 => conv1_dout_net_x0,
      in2 => conv2_dout_net_x0,
      in3 => conv3_dout_net_x0,
      in4 => conv4_dout_net_x0,
      bus_out => concatenate_y_net_x1
    );

  conv1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x99,
      clk => clk_1_sg_x99,
      clr => '0',
      din => reinterpret4_output_port_net_x0,
      en => "1",
      dout => conv1_dout_net_x0
    );

  conv2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x99,
      clk => clk_1_sg_x99,
      clr => '0',
      din => reinterpret3_output_port_net_x0,
      en => "1",
      dout => conv2_dout_net_x0
    );

  conv3: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x99,
      clk => clk_1_sg_x99,
      clr => '0',
      din => reinterpret2_output_port_net_x0,
      en => "1",
      dout => conv3_dout_net_x0
    );

  conv4: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 17,
      din_width => 20,
      dout_arith => 2,
      dout_bin_pt => 18,
      dout_width => 21,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x99,
      clk => clk_1_sg_x99,
      clr => '0',
      din => reinterpret1_output_port_net_x0,
      en => "1",
      dout => conv4_dout_net_x0
    );

  debus_fe21c1b916: entity work.debus_entity_fe21c1b916
    port map (
      bus_in => concat_y_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_norm1/conv1"

entity conv1_entity_75f0e5795b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(19 downto 0); 
    out_x0: out std_logic_vector(20 downto 0)
  );
end conv1_entity_75f0e5795b;

architecture structural of conv1_entity_75f0e5795b is
  signal adder_s_net_x4: std_logic_vector(20 downto 0);
  signal almost_half_op_net: std_logic_vector(18 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x100: std_logic;
  signal clk_1_sg_x100: std_logic;
  signal concat_y_net: std_logic_vector(20 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(20 downto 0);
  signal force2_output_port_net: std_logic_vector(18 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(19 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x100 <= ce_1;
  clk_1_sg_x100 <= clk_1;
  reinterpret4_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x4;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 19,
      a_width => 21,
      b_arith => xlUnsigned,
      b_bin_pt => 19,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 22,
      core_name0 => "addsb_11_0_c055560701350b3e",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 22,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 18,
      s_width => 21
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x100,
      clk => clk_1_sg_x100,
      clr => '0',
      en => "1",
      s => adder_s_net_x4
    );

  almost_half: entity work.constant_b366689086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 20,
      y_width => 1
    )
    port map (
      x => reinterpret4_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_c615d93998
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_d357e69fa3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_d2180c9169
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_4a8cbc85ce
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret4_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_b1e9d7c303
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_norm1"

entity bus_norm1_entity_cc02258db8 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(83 downto 0)
  );
end bus_norm1_entity_cc02258db8;

architecture structural of bus_norm1_entity_cc02258db8 is
  signal adder_s_net_x4: std_logic_vector(20 downto 0);
  signal adder_s_net_x5: std_logic_vector(20 downto 0);
  signal adder_s_net_x6: std_logic_vector(20 downto 0);
  signal adder_s_net_x7: std_logic_vector(20 downto 0);
  signal ce_1_sg_x104: std_logic;
  signal clk_1_sg_x104: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(19 downto 0);

begin
  ce_1_sg_x104 <= ce_1;
  clk_1_sg_x104 <= clk_1;
  concatenate_y_net_x2 <= din;
  dout <= concatenate_y_net_x3;

  bussify_2e70185336: entity work.bussify_entity_83bee71966
    port map (
      in1 => adder_s_net_x4,
      in2 => adder_s_net_x5,
      in3 => adder_s_net_x6,
      in4 => adder_s_net_x7,
      bus_out => concatenate_y_net_x3
    );

  conv1_75f0e5795b: entity work.conv1_entity_75f0e5795b
    port map (
      ce_1 => ce_1_sg_x104,
      clk_1 => clk_1_sg_x104,
      in_x0 => reinterpret4_output_port_net_x1,
      out_x0 => adder_s_net_x4
    );

  conv2_c4ef7f773d: entity work.conv1_entity_75f0e5795b
    port map (
      ce_1 => ce_1_sg_x104,
      clk_1 => clk_1_sg_x104,
      in_x0 => reinterpret3_output_port_net_x1,
      out_x0 => adder_s_net_x5
    );

  conv3_d40d6825c2: entity work.conv1_entity_75f0e5795b
    port map (
      ce_1 => ce_1_sg_x104,
      clk_1 => clk_1_sg_x104,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x6
    );

  conv4_f8c41adab0: entity work.conv1_entity_75f0e5795b
    port map (
      ce_1 => ce_1_sg_x104,
      clk_1 => clk_1_sg_x104,
      in_x0 => reinterpret1_output_port_net_x1,
      out_x0 => adder_s_net_x7
    );

  debus_661a1cbfb6: entity work.debus_entity_5abef6bede
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_scale"

entity bus_scale_entity_5b3b5027bd is
  port (
    din: in std_logic_vector(79 downto 0); 
    dout: out std_logic_vector(79 downto 0)
  );
end bus_scale_entity_5b3b5027bd;

architecture structural of bus_scale_entity_5b3b5027bd is
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(19 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(19 downto 0);
  signal scale1_op_net_x0: std_logic_vector(19 downto 0);
  signal scale2_op_net_x0: std_logic_vector(19 downto 0);
  signal scale3_op_net_x0: std_logic_vector(19 downto 0);
  signal scale4_op_net_x0: std_logic_vector(19 downto 0);

begin
  concat_y_net_x3 <= din;
  dout <= concatenate_y_net_x4;

  bussify_d65e371524: entity work.bussify_entity_c32f93b775
    port map (
      in1 => scale1_op_net_x0,
      in2 => scale2_op_net_x0,
      in3 => scale3_op_net_x0,
      in4 => scale4_op_net_x0,
      bus_out => concatenate_y_net_x4
    );

  debus_3211bd7379: entity work.debus_entity_fe21c1b916
    port map (
      bus_in => concat_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  scale1: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret4_output_port_net_x0,
      op => scale1_op_net_x0
    );

  scale2: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret3_output_port_net_x0,
      op => scale2_op_net_x0
    );

  scale3: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret2_output_port_net_x0,
      op => scale3_op_net_x0
    );

  scale4: entity work.scale_97239b8ed2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      ip => reinterpret1_output_port_net_x0,
      op => scale4_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/bus_sub"

entity bus_sub_entity_041fbb1680 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(37 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dout: out std_logic_vector(39 downto 0)
  );
end bus_sub_entity_041fbb1680;

architecture structural of bus_sub_entity_041fbb1680 is
  signal addsub1_s_net_x0: std_logic_vector(19 downto 0);
  signal addsub2_s_net_x0: std_logic_vector(19 downto 0);
  signal ce_1_sg_x105: std_logic;
  signal clk_1_sg_x105: std_logic;
  signal concatenate_y_net_x4: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(39 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(18 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(18 downto 0);

begin
  reinterpret1_output_port_net_x5 <= a;
  concatenate_y_net_x4 <= b;
  ce_1_sg_x105 <= ce_1;
  clk_1_sg_x105 <= clk_1;
  dout <= concatenate_y_net_x5;

  a_debus_682093e7bc: entity work.a_debus_entity_e8ca01a28d
    port map (
      bus_in => reinterpret1_output_port_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x0
    );

  addsub1: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_a0497faccc62b6b2",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x105,
      clk => clk_1_sg_x105,
      clr => '0',
      en => "1",
      s => addsub1_s_net_x0
    );

  addsub2: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 17,
      a_width => 18,
      b_arith => xlSigned,
      b_bin_pt => 17,
      b_width => 19,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 20,
      core_name0 => "addsb_11_0_a0497faccc62b6b2",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 20,
      latency => 2,
      overflow => 2,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 20
    )
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret1_output_port_net_x1,
      ce => ce_1_sg_x105,
      clk => clk_1_sg_x105,
      clr => '0',
      en => "1",
      s => addsub2_s_net_x0
    );

  b_debus_e9034d57c1: entity work.b_debus_entity_97187af928
    port map (
      bus_in => concatenate_y_net_x4,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  op_bussify_c96c03eb4c: entity work.op_bussify_entity_cf1986e0b4
    port map (
      in1 => addsub1_s_net_x0,
      in2 => addsub2_s_net_x0,
      bus_out => concatenate_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/mux/d_bussify"

entity d_bussify_entity_66e7d11cd7 is
  port (
    in1: in std_logic_vector(20 downto 0); 
    in2: in std_logic_vector(20 downto 0); 
    in3: in std_logic_vector(20 downto 0); 
    in4: in std_logic_vector(20 downto 0); 
    bus_out: out std_logic_vector(83 downto 0)
  );
end d_bussify_entity_66e7d11cd7;

architecture structural of d_bussify_entity_66e7d11cd7 is
  signal concatenate_y_net_x4: std_logic_vector(83 downto 0);
  signal mux0_y_net_x0: std_logic_vector(20 downto 0);
  signal mux1_y_net_x0: std_logic_vector(20 downto 0);
  signal mux2_y_net_x0: std_logic_vector(20 downto 0);
  signal mux3_y_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(20 downto 0);

begin
  mux0_y_net_x0 <= in1;
  mux1_y_net_x0 <= in2;
  mux2_y_net_x0 <= in3;
  mux3_y_net_x0 <= in4;
  bus_out <= concatenate_y_net_x4;

  concatenate: entity work.concat_356a264444
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x4
    );

  reinterpret1: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux0_y_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux1_y_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux2_y_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux3_y_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/mux/expand0"

entity expand0_entity_bede1f0eab is
  port (
    bus_in: in std_logic_vector(83 downto 0); 
    lsb_out1: out std_logic_vector(20 downto 0); 
    msb_out4: out std_logic_vector(20 downto 0); 
    out2: out std_logic_vector(20 downto 0); 
    out3: out std_logic_vector(20 downto 0)
  );
end expand0_entity_bede1f0eab;

architecture structural of expand0_entity_bede1f0eab is
  signal concatenate_y_net_x2: std_logic_vector(83 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(20 downto 0);
  signal slice1_y_net: std_logic_vector(20 downto 0);
  signal slice2_y_net: std_logic_vector(20 downto 0);
  signal slice3_y_net: std_logic_vector(20 downto 0);
  signal slice4_y_net: std_logic_vector(20 downto 0);

begin
  concatenate_y_net_x2 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_299ca43e25
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 20,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 21,
      new_msb => 41,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 42,
      new_msb => 62,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 63,
      new_msb => 83,
      x_width => 84,
      y_width => 21
    )
    port map (
      x => concatenate_y_net_x2,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/mux"

entity mux_entity_2a2e20cd83 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d0: in std_logic_vector(83 downto 0); 
    d1: in std_logic_vector(83 downto 0); 
    sel: in std_logic_vector(3 downto 0); 
    out_x0: out std_logic_vector(83 downto 0)
  );
end mux_entity_2a2e20cd83;

architecture structural of mux_entity_2a2e20cd83 is
  signal ce_1_sg_x106: std_logic;
  signal clk_1_sg_x106: std_logic;
  signal concatenate_y_net_x6: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(83 downto 0);
  signal mux0_y_net_x0: std_logic_vector(20 downto 0);
  signal mux1_y_net_x0: std_logic_vector(20 downto 0);
  signal mux2_y_net_x0: std_logic_vector(20 downto 0);
  signal mux3_y_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(20 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(20 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic;
  signal reinterpret3_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(20 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic;
  signal reinterpret4_output_port_net_x0: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(20 downto 0);
  signal reinterpret4_output_port_net_x2: std_logic;

begin
  ce_1_sg_x106 <= ce_1;
  clk_1_sg_x106 <= clk_1;
  concatenate_y_net_x6 <= d0;
  concatenate_y_net_x7 <= d1;
  concatenate_y_net_x8 <= sel;
  out_x0 <= concatenate_y_net_x9;

  d_bussify_66e7d11cd7: entity work.d_bussify_entity_66e7d11cd7
    port map (
      in1 => mux0_y_net_x0,
      in2 => mux1_y_net_x0,
      in3 => mux2_y_net_x0,
      in4 => mux3_y_net_x0,
      bus_out => concatenate_y_net_x9
    );

  expand0_bede1f0eab: entity work.expand0_entity_bede1f0eab
    port map (
      bus_in => concatenate_y_net_x6,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  expand1_89b5d0e2c9: entity work.expand0_entity_bede1f0eab
    port map (
      bus_in => concatenate_y_net_x7,
      lsb_out1 => reinterpret1_output_port_net_x1,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

  mux0: entity work.mux_46aae2a33a
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      d0 => reinterpret4_output_port_net_x0,
      d1 => reinterpret4_output_port_net_x1,
      sel(0) => reinterpret4_output_port_net_x2,
      y => mux0_y_net_x0
    );

  mux1: entity work.mux_46aae2a33a
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      d0 => reinterpret3_output_port_net_x0,
      d1 => reinterpret3_output_port_net_x1,
      sel(0) => reinterpret3_output_port_net_x2,
      y => mux1_y_net_x0
    );

  mux2: entity work.mux_46aae2a33a
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      d0 => reinterpret2_output_port_net_x0,
      d1 => reinterpret2_output_port_net_x1,
      sel(0) => reinterpret2_output_port_net_x2,
      y => mux2_y_net_x0
    );

  mux3: entity work.mux_46aae2a33a
    port map (
      ce => ce_1_sg_x106,
      clk => clk_1_sg_x106,
      clr => '0',
      d0 => reinterpret1_output_port_net_x0,
      d1 => reinterpret1_output_port_net_x1,
      sel(0) => reinterpret1_output_port_net_x2,
      y => mux3_y_net_x0
    );

  sel_expand_23a6ff5fd7: entity work.sel_expand_entity_41b2560930
    port map (
      bus_in => concatenate_y_net_x8,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out4 => reinterpret4_output_port_net_x2,
      out2 => reinterpret2_output_port_net_x2,
      out3 => reinterpret3_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert/conv1"

entity conv1_entity_d275b9050a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(36 downto 0); 
    out_x0: out std_logic_vector(18 downto 0)
  );
end conv1_entity_d275b9050a;

architecture structural of conv1_entity_d275b9050a is
  signal adder_s_net_x2: std_logic_vector(18 downto 0);
  signal almost_half_op_net: std_logic_vector(34 downto 0);
  signal bit_y_net: std_logic;
  signal ce_1_sg_x108: std_logic;
  signal clk_1_sg_x108: std_logic;
  signal concat_y_net: std_logic_vector(37 downto 0);
  signal constant_op_net: std_logic;
  signal force1_output_port_net: std_logic_vector(37 downto 0);
  signal force2_output_port_net: std_logic_vector(34 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(36 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(36 downto 0);
  signal tweak_op_y_net: std_logic;

begin
  ce_1_sg_x108 <= ce_1;
  clk_1_sg_x108 <= clk_1;
  reinterpret2_output_port_net_x0 <= in_x0;
  out_x0 <= adder_s_net_x2;

  adder: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 35,
      a_width => 38,
      b_arith => xlUnsigned,
      b_bin_pt => 35,
      b_width => 35,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 39,
      core_name0 => "addsb_11_0_6e641a09b813308f",
      extra_registers => 1,
      full_s_arith => 2,
      full_s_width => 39,
      latency => 2,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 17,
      s_width => 19
    )
    port map (
      a => force1_output_port_net,
      b => force2_output_port_net,
      ce => ce_1_sg_x108,
      clk => clk_1_sg_x108,
      clr => '0',
      en => "1",
      s => adder_s_net_x2
    );

  almost_half: entity work.constant_2da6af93c2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => almost_half_op_net
    );

  bit: entity work.xlslice
    generic map (
      new_lsb => 17,
      new_msb => 17,
      x_width => 37,
      y_width => 1
    )
    port map (
      x => reinterpret2_output_port_net_x0,
      y(0) => bit_y_net
    );

  concat: entity work.concat_83820b2faf
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1(0) => tweak_op_y_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  force1: entity work.reinterpret_620dd01637
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => force1_output_port_net
    );

  force2: entity work.reinterpret_ec14c62a89
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => almost_half_op_net,
      output_port => force2_output_port_net
    );

  reinterpret: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret2_output_port_net_x0,
      output_port => reinterpret_output_port_net
    );

  tweak_op: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => bit_y_net,
      d1(0) => constant_op_net,
      y(0) => tweak_op_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert/debus"

entity debus_entity_af63b30568 is
  port (
    bus_in: in std_logic_vector(73 downto 0); 
    lsb_out1: out std_logic_vector(36 downto 0); 
    msb_out2: out std_logic_vector(36 downto 0)
  );
end debus_entity_af63b30568;

architecture structural of debus_entity_af63b30568 is
  signal reinterpret1_output_port_net_x1: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(36 downto 0);
  signal slice1_y_net: std_logic_vector(36 downto 0);
  signal slice2_y_net: std_logic_vector(36 downto 0);

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x2;
  msb_out2 <= reinterpret2_output_port_net_x1;

  reinterpret1: entity work.reinterpret_5b4829fb41
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  reinterpret2: entity work.reinterpret_5b4829fb41
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 36,
      x_width => 74,
      y_width => 37
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 37,
      new_msb => 73,
      x_width => 74,
      y_width => 37
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_convert"

entity bus_convert_entity_e5fd0829de is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(73 downto 0); 
    misci: in std_logic_vector(36 downto 0); 
    dout: out std_logic_vector(37 downto 0); 
    misco: out std_logic_vector(36 downto 0)
  );
end bus_convert_entity_e5fd0829de;

architecture structural of bus_convert_entity_e5fd0829de is
  signal adder_s_net_x2: std_logic_vector(18 downto 0);
  signal adder_s_net_x3: std_logic_vector(18 downto 0);
  signal ce_1_sg_x110: std_logic;
  signal clk_1_sg_x110: std_logic;
  signal concatenate_y_net_x6: std_logic_vector(37 downto 0);
  signal dmisc_q_net_x1: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(73 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(36 downto 0);

begin
  ce_1_sg_x110 <= ce_1;
  clk_1_sg_x110 <= clk_1;
  reinterpret1_output_port_net_x3 <= din;
  dmisc_q_net_x1 <= misci;
  dout <= concatenate_y_net_x6;
  misco <= dmisc_q_net_x2;

  bussify_a0ef8580a2: entity work.op_bussify_entity_a6d4bedd3c
    port map (
      in1 => adder_s_net_x2,
      in2 => adder_s_net_x3,
      bus_out => concatenate_y_net_x6
    );

  conv1_d275b9050a: entity work.conv1_entity_d275b9050a
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      in_x0 => reinterpret2_output_port_net_x1,
      out_x0 => adder_s_net_x2
    );

  conv2_ad83469104: entity work.conv1_entity_d275b9050a
    port map (
      ce_1 => ce_1_sg_x110,
      clk_1 => clk_1_sg_x110,
      in_x0 => reinterpret1_output_port_net_x2,
      out_x0 => adder_s_net_x3
    );

  debus_af63b30568: entity work.debus_entity_af63b30568
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x2,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  dmisc: entity work.delay_8e134646d3
    port map (
      ce => ce_1_sg_x110,
      clk => clk_1_sg_x110,
      clr => '0',
      d => dmisc_q_net_x1,
      q => dmisc_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_create"

entity bus_create_entity_1ff518d55f is
  port (
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic; 
    in3: in std_logic_vector(35 downto 0); 
    bus_out: out std_logic_vector(72 downto 0)
  );
end bus_create_entity_1ff518d55f;

architecture structural of bus_create_entity_1ff518d55f is
  signal concatenate_y_net_x0: std_logic_vector(72 downto 0);
  signal dmux0_q_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x0: std_logic;
  signal reinterpret1_output_port_net: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net: std_logic;
  signal reinterpret3_output_port_net: std_logic_vector(35 downto 0);

begin
  dmux0_q_net_x0 <= in1;
  mux_y_net_x0 <= in2;
  reinterpret1_output_port_net_x1 <= in3;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_b28df1ab2e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1(0) => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => dmux0_q_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_112d91c147
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port(0) => mux_y_net_x0,
      output_port(0) => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => reinterpret1_output_port_net_x1,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_expand"

entity bus_expand_entity_56cf888bad is
  port (
    bus_in: in std_logic_vector(72 downto 0); 
    lsb_out1: out std_logic_vector(36 downto 0); 
    msb_out2: out std_logic_vector(35 downto 0)
  );
end bus_expand_entity_56cf888bad;

architecture structural of bus_expand_entity_56cf888bad is
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(36 downto 0);
  signal slice2_y_net: std_logic_vector(35 downto 0);

begin
  delay1_q_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out2 <= reinterpret2_output_port_net_x0;

  reinterpret1: entity work.reinterpret_892b735f0d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 36,
      x_width => 73,
      y_width => 37
    )
    port map (
      x => delay1_q_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 37,
      new_msb => 72,
      x_width => 73,
      y_width => 36
    )
    port map (
      x => delay1_q_net_x0,
      y => slice2_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_expand1"

entity bus_expand1_entity_bcd05ee4e4 is
  port (
    bus_in: in std_logic_vector(36 downto 0); 
    lsb_out1: out std_logic_vector(35 downto 0); 
    msb_out2: out std_logic
  );
end bus_expand1_entity_bcd05ee4e4;

architecture structural of bus_expand1_entity_bcd05ee4e4 is
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice1_y_net: std_logic_vector(35 downto 0);
  signal slice2_y_net_x0: std_logic;

begin
  dmisc_q_net_x3 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x6;
  msb_out2 <= slice2_y_net_x0;

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x6
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 35,
      x_width => 37,
      y_width => 36
    )
    port map (
      x => dmisc_q_net_x3,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 36,
      x_width => 37,
      y_width => 1
    )
    port map (
      x => dmisc_q_net_x3,
      y(0) => slice2_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/a*b_bussify"

entity a_b_bussify_entity_5f7d61d0c0 is
  port (
    in1: in std_logic_vector(73 downto 0); 
    bus_out: out std_logic_vector(73 downto 0)
  );
end a_b_bussify_entity_5f7d61d0c0;

architecture structural of a_b_bussify_entity_5f7d61d0c0 is
  signal concat_y_net_x0: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(73 downto 0);

begin
  concat_y_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x4;

  reinterpret1: entity work.reinterpret_efdf1c3890
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net_x0,
      output_port => reinterpret1_output_port_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/a_expand"

entity a_expand_entity_69cb316c5d is
  port (
    bus_in: in std_logic_vector(71 downto 0); 
    lsb_out1: out std_logic_vector(17 downto 0); 
    msb_out4: out std_logic_vector(17 downto 0); 
    out2: out std_logic_vector(17 downto 0); 
    out3: out std_logic_vector(17 downto 0)
  );
end a_expand_entity_69cb316c5d;

architecture structural of a_expand_entity_69cb316c5d is
  signal concatenate_y_net_x0: std_logic_vector(71 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(17 downto 0);
  signal slice1_y_net: std_logic_vector(17 downto 0);
  signal slice2_y_net: std_logic_vector(17 downto 0);
  signal slice3_y_net: std_logic_vector(17 downto 0);
  signal slice4_y_net: std_logic_vector(17 downto 0);

begin
  concatenate_y_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 36,
      new_msb => 53,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 54,
      new_msb => 71,
      x_width => 72,
      y_width => 18
    )
    port map (
      x => concatenate_y_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/a_replicate/bussify"

entity bussify_entity_a3555039c4 is
  port (
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    bus_out: out std_logic_vector(71 downto 0)
  );
end bussify_entity_a3555039c4;

architecture structural of bussify_entity_a3555039c4 is
  signal concatenate_y_net_x1: std_logic_vector(71 downto 0);
  signal din0_0_q_net_x0: std_logic_vector(35 downto 0);
  signal din0_1_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(35 downto 0);

begin
  din0_0_q_net_x0 <= in1;
  din0_1_q_net_x0 <= in2;
  bus_out <= concatenate_y_net_x1;

  concatenate: entity work.concat_c3ccc04d1a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      y => concatenate_y_net_x1
    );

  reinterpret1: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din0_0_q_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_86b044698f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din0_1_q_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/a_replicate"

entity a_replicate_entity_aa69b6fc2b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(35 downto 0); 
    out_x0: out std_logic_vector(71 downto 0)
  );
end a_replicate_entity_aa69b6fc2b;

architecture structural of a_replicate_entity_aa69b6fc2b is
  signal ce_1_sg_x111: std_logic;
  signal clk_1_sg_x111: std_logic;
  signal concatenate_y_net_x2: std_logic_vector(71 downto 0);
  signal din0_0_q_net_x0: std_logic_vector(35 downto 0);
  signal din0_1_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x111 <= ce_1;
  clk_1_sg_x111 <= clk_1;
  reinterpret1_output_port_net_x3 <= in_x0;
  out_x0 <= concatenate_y_net_x2;

  bussify_a3555039c4: entity work.bussify_entity_a3555039c4
    port map (
      in1 => din0_0_q_net_x0,
      in2 => din0_1_q_net_x0,
      bus_out => concatenate_y_net_x2
    );

  din0_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 36
    )
    port map (
      ce => ce_1_sg_x111,
      clk => clk_1_sg_x111,
      d => reinterpret1_output_port_net_x3,
      en => '1',
      rst => '1',
      q => din0_0_q_net_x0
    );

  din0_1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 36
    )
    port map (
      ce => ce_1_sg_x111,
      clk => clk_1_sg_x111,
      d => reinterpret1_output_port_net_x3,
      en => '1',
      rst => '1',
      q => din0_1_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1/ri_to_c"

entity ri_to_c_entity_8ac70ac307 is
  port (
    im: in std_logic_vector(36 downto 0); 
    re: in std_logic_vector(36 downto 0); 
    c: out std_logic_vector(73 downto 0)
  );
end ri_to_c_entity_8ac70ac307;

architecture structural of ri_to_c_entity_8ac70ac307 is
  signal concat_y_net_x1: std_logic_vector(73 downto 0);
  signal convert_im_dout_net_x0: std_logic_vector(36 downto 0);
  signal convert_re_dout_net_x0: std_logic_vector(36 downto 0);
  signal force_im_output_port_net: std_logic_vector(36 downto 0);
  signal force_re_output_port_net: std_logic_vector(36 downto 0);

begin
  convert_im_dout_net_x0 <= im;
  convert_re_dout_net_x0 <= re;
  c <= concat_y_net_x1;

  concat: entity work.concat_56d57d2c92
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x1
    );

  force_im: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_im_dout_net_x0,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_db4c53ade5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_re_dout_net_x0,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/mult1"

entity mult1_entity_72a01a3ec3 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    ab: out std_logic_vector(73 downto 0)
  );
end mult1_entity_72a01a3ec3;

architecture structural of mult1_entity_72a01a3ec3 is
  signal addsub_im_s_net: std_logic_vector(36 downto 0);
  signal addsub_re_s_net: std_logic_vector(36 downto 0);
  signal ce_1_sg_x113: std_logic;
  signal clk_1_sg_x113: std_logic;
  signal concat_y_net_x2: std_logic_vector(73 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(71 downto 0);
  signal convert_im_dout_net_x0: std_logic_vector(36 downto 0);
  signal convert_re_dout_net_x0: std_logic_vector(36 downto 0);
  signal imim_p_net: std_logic_vector(35 downto 0);
  signal imre_p_net: std_logic_vector(35 downto 0);
  signal reim_p_net: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(17 downto 0);
  signal rere_p_net: std_logic_vector(35 downto 0);

begin
  reinterpret1_output_port_net_x6 <= a;
  reinterpret1_output_port_net_x7 <= b;
  ce_1_sg_x113 <= ce_1;
  clk_1_sg_x113 <= clk_1;
  ab <= concat_y_net_x2;

  a_expand_69cb316c5d: entity work.a_expand_entity_69cb316c5d
    port map (
      bus_in => concatenate_y_net_x2,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  a_replicate_aa69b6fc2b: entity work.a_replicate_entity_aa69b6fc2b
    port map (
      ce_1 => ce_1_sg_x113,
      clk_1 => clk_1_sg_x113,
      in_x0 => reinterpret1_output_port_net_x6,
      out_x0 => concatenate_y_net_x2
    );

  addsub_im: entity work.addsub_4ded11ba54
    port map (
      a => imre_p_net,
      b => reim_p_net,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      s => addsub_im_s_net
    );

  addsub_re: entity work.addsub_8dd4a43ef5
    port map (
      a => rere_p_net,
      b => imim_p_net,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      s => addsub_re_s_net
    );

  b_expand_00682737c0: entity work.a_expand_entity_69cb316c5d
    port map (
      bus_in => concatenate_y_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out4 => reinterpret4_output_port_net_x1,
      out2 => reinterpret2_output_port_net_x1,
      out3 => reinterpret3_output_port_net_x1
    );

  b_replicate_595c449808: entity work.a_replicate_entity_aa69b6fc2b
    port map (
      ce_1 => ce_1_sg_x113,
      clk_1 => clk_1_sg_x113,
      in_x0 => reinterpret1_output_port_net_x7,
      out_x0 => concatenate_y_net_x3
    );

  convert_im: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 34,
      din_width => 37,
      dout_arith => 2,
      dout_bin_pt => 34,
      dout_width => 37,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      din => addsub_im_s_net,
      en => "1",
      dout => convert_im_dout_net_x0
    );

  convert_re: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 34,
      din_width => 37,
      dout_arith => 2,
      dout_bin_pt => 34,
      dout_width => 37,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      din => addsub_re_s_net,
      en => "1",
      dout => convert_re_dout_net_x0
    );

  imim: entity work.mult_f295e5f0f2
    port map (
      a => reinterpret3_output_port_net_x0,
      b => reinterpret3_output_port_net_x1,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      p => imim_p_net
    );

  imre: entity work.mult_f295e5f0f2
    port map (
      a => reinterpret1_output_port_net_x0,
      b => reinterpret2_output_port_net_x1,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      p => imre_p_net
    );

  reim: entity work.mult_f295e5f0f2
    port map (
      a => reinterpret2_output_port_net_x0,
      b => reinterpret1_output_port_net_x5,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      p => reim_p_net
    );

  rere: entity work.mult_f295e5f0f2
    port map (
      a => reinterpret4_output_port_net_x0,
      b => reinterpret4_output_port_net_x1,
      ce => ce_1_sg_x113,
      clk => clk_1_sg_x113,
      clr => '0',
      p => rere_p_net
    );

  ri_to_c_8ac70ac307: entity work.ri_to_c_entity_8ac70ac307
    port map (
      im => convert_im_dout_net_x0,
      re => convert_re_dout_net_x0,
      c => concat_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult/repa"

entity repa_entity_d74ee50680 is
  port (
    in_x0: in std_logic_vector(35 downto 0); 
    out_x0: out std_logic_vector(35 downto 0)
  );
end repa_entity_d74ee50680;

architecture structural of repa_entity_d74ee50680 is
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);

begin
  concat_y_net_x1 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x3;

  bussify_63e56c0409: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => concat_y_net_x1,
      bus_out => reinterpret1_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/bus_mult"

entity bus_mult_entity_b0541e7d96 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(36 downto 0); 
    a_b: out std_logic_vector(73 downto 0); 
    misco: out std_logic_vector(36 downto 0)
  );
end bus_mult_entity_b0541e7d96;

architecture structural of bus_mult_entity_b0541e7d96 is
  signal ce_1_sg_x114: std_logic;
  signal clk_1_sg_x114: std_logic;
  signal concat_y_net_x2: std_logic_vector(73 downto 0);
  signal concat_y_net_x3: std_logic_vector(35 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);

begin
  concat_y_net_x3 <= a;
  reinterpret2_output_port_net_x3 <= b;
  ce_1_sg_x114 <= ce_1;
  clk_1_sg_x114 <= clk_1;
  reinterpret1_output_port_net_x9 <= misci;
  a_b <= reinterpret1_output_port_net_x10;
  misco <= dmisc_q_net_x2;

  a_b_bussify_5f7d61d0c0: entity work.a_b_bussify_entity_5f7d61d0c0
    port map (
      in1 => concat_y_net_x2,
      bus_out => reinterpret1_output_port_net_x10
    );

  a_debus_2a36773c9a: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x6
    );

  b_debus_3d6035e944: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x8,
      msb_lsb_out1 => reinterpret1_output_port_net_x7
    );

  dmisc: entity work.delay_2d0f74b2c1
    port map (
      ce => ce_1_sg_x114,
      clk => clk_1_sg_x114,
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => dmisc_q_net_x2
    );

  mult1_72a01a3ec3: entity work.mult1_entity_72a01a3ec3
    port map (
      a => reinterpret1_output_port_net_x6,
      b => reinterpret1_output_port_net_x7,
      ce_1 => ce_1_sg_x114,
      clk_1 => clk_1_sg_x114,
      ab => concat_y_net_x2
    );

  repa_d74ee50680: entity work.repa_entity_d74ee50680
    port map (
      in_x0 => concat_y_net_x3,
      out_x0 => reinterpret1_output_port_net_x3
    );

  repb_c759917e7d: entity work.repa_entity_d74ee50680
    port map (
      in_x0 => reinterpret2_output_port_net_x3,
      out_x0 => reinterpret1_output_port_net_x8
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_f05b79004d is
  port (
    in_x0: in std_logic_vector(8 downto 0); 
    out_x0: out std_logic_vector(8 downto 0)
  );
end bit_reverse_entity_f05b79004d;

architecture structural of bit_reverse_entity_f05b79004d is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(8 downto 0);
  signal slice_y_net_x0: std_logic_vector(8 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  concat: entity work.concat_0cc72cd991
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_6677c7a36d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(8 downto 0); 
    add: out std_logic_vector(8 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_6677c7a36d;

architecture structural of add_convert0_entity_6677c7a36d is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(8 downto 0);
  signal ce_1_sg_x115: std_logic;
  signal clk_1_sg_x115: std_logic;
  signal concat_y_net: std_logic_vector(9 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal delay13_q_net: std_logic_vector(8 downto 0);
  signal delay14_q_net: std_logic_vector(8 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(9 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(7 downto 0);
  signal new_add_y_net: std_logic_vector(8 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x115 <= ce_1;
  clk_1_sg_x115 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x115,
      clk => clk_1_sg_x115,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_7eef56098d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 9,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 9,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x115,
      clk => clk_1_sg_x115,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_6104cbef7a
    port map (
      ce => ce_1_sg_x115,
      clk => clk_1_sg_x115,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_09771002d6
    port map (
      ce => ce_1_sg_x115,
      clk => clk_1_sg_x115,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x115,
      clk => clk_1_sg_x115,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9779a5cf83
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 10,
      y_width => 8
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 10,
      y_width => 9
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 9,
      x_width => 10,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_9b7575767f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(8 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_9b7575767f;

architecture structural of add_convert1_entity_9b7575767f is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x116: std_logic;
  signal clk_1_sg_x116: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(9 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x116 <= ce_1;
  clk_1_sg_x116 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x116,
      clk => clk_1_sg_x116,
      clr => '0',
      s => addsub5_s_net
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x116,
      clk => clk_1_sg_x116,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x116,
      clk => clk_1_sg_x116,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9779a5cf83
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 9,
      x_width => 10,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/c_to_ri"

entity c_to_ri_entity_ef07e318f3 is
  port (
    c: in std_logic_vector(35 downto 0); 
    im: out std_logic_vector(17 downto 0); 
    re: out std_logic_vector(17 downto 0)
  );
end c_to_ri_entity_ef07e318f3;

architecture structural of c_to_ri_entity_ef07e318f3 is
  signal force_im_output_port_net_x0: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x0: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);
  signal slice_im_y_net: std_logic_vector(17 downto 0);
  signal slice_re_y_net: std_logic_vector(17 downto 0);

begin
  rom_data_net_x0 <= c;
  im <= force_im_output_port_net_x0;
  re <= force_re_output_port_net_x0;

  force_im: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_im_y_net,
      output_port => force_im_output_port_net_x0
    );

  force_re: entity work.reinterpret_9a0fa0f632
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_re_y_net,
      output_port => force_re_output_port_net_x0
    );

  slice_im: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 17,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => rom_data_net_x0,
      y => slice_im_y_net
    );

  slice_re: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 35,
      x_width => 36,
      y_width => 18
    )
    port map (
      x => rom_data_net_x0,
      y => slice_re_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/invert0"

entity invert0_entity_00bc692256 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(17 downto 0); 
    negate_x0: in std_logic; 
    out_x0: out std_logic_vector(17 downto 0)
  );
end invert0_entity_00bc692256;

architecture structural of invert0_entity_00bc692256 is
  signal ce_1_sg_x117: std_logic;
  signal clk_1_sg_x117: std_logic;
  signal delay10_q_net_x0: std_logic;
  signal delay20_q_net: std_logic_vector(17 downto 0);
  signal delay21_q_net: std_logic;
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x0: std_logic_vector(17 downto 0);
  signal negate_op_net: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x117 <= ce_1;
  clk_1_sg_x117 <= clk_1;
  force_re_output_port_net_x1 <= in_x0;
  delay10_q_net_x0 <= negate_x0;
  out_x0 <= mux_y_net_x0;

  delay20: entity work.delay_b6092ad150
    port map (
      ce => ce_1_sg_x117,
      clk => clk_1_sg_x117,
      clr => '0',
      d => force_re_output_port_net_x1,
      q => delay20_q_net
    );

  delay21: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x117,
      clk => clk_1_sg_x117,
      clr => '0',
      d(0) => delay10_q_net_x0,
      q(0) => delay21_q_net
    );

  mux: entity work.mux_1896e7760c
    port map (
      ce => ce_1_sg_x117,
      clk => clk_1_sg_x117,
      clr => '0',
      d0 => delay20_q_net,
      d1 => negate_op_net,
      sel(0) => delay21_q_net,
      y => mux_y_net_x0
    );

  negate: entity work.negate_206b7f76d8
    port map (
      ce => ce_1_sg_x117,
      clk => clk_1_sg_x117,
      clr => '0',
      ip => force_re_output_port_net_x1,
      op => negate_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin/invert1"

entity invert1_entity_17dc85599c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(17 downto 0); 
    misci: in std_logic_vector(72 downto 0); 
    negate_x0: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    out_x0: out std_logic_vector(17 downto 0)
  );
end invert1_entity_17dc85599c;

architecture structural of invert1_entity_17dc85599c is
  signal ce_1_sg_x118: std_logic;
  signal clk_1_sg_x118: std_logic;
  signal delay1_q_net_x1: std_logic_vector(72 downto 0);
  signal delay20_q_net: std_logic_vector(17 downto 0);
  signal delay21_q_net: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x0: std_logic_vector(17 downto 0);
  signal negate_op_net: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x118 <= ce_1;
  clk_1_sg_x118 <= clk_1;
  force_im_output_port_net_x1 <= in_x0;
  delay_q_net_x0 <= misci;
  delay8_q_net_x0 <= negate_x0;
  misco <= delay1_q_net_x1;
  out_x0 <= mux_y_net_x0;

  delay1: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x118,
      clk => clk_1_sg_x118,
      clr => '0',
      d => delay_q_net_x0,
      q => delay1_q_net_x1
    );

  delay20: entity work.delay_b6092ad150
    port map (
      ce => ce_1_sg_x118,
      clk => clk_1_sg_x118,
      clr => '0',
      d => force_im_output_port_net_x1,
      q => delay20_q_net
    );

  delay21: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x118,
      clk => clk_1_sg_x118,
      clr => '0',
      d(0) => delay8_q_net_x0,
      q(0) => delay21_q_net
    );

  mux: entity work.mux_1896e7760c
    port map (
      ce => ce_1_sg_x118,
      clk => clk_1_sg_x118,
      clr => '0',
      d0 => delay20_q_net,
      d1 => negate_op_net,
      sel(0) => delay21_q_net,
      y => mux_y_net_x0
    );

  negate: entity work.negate_206b7f76d8
    port map (
      ce => ce_1_sg_x118,
      clk => clk_1_sg_x118,
      clr => '0',
      ip => force_im_output_port_net_x1,
      op => negate_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_8c6d36a3ce is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(8 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_8c6d36a3ce;

architecture structural of cosin_entity_8c6d36a3ce is
  signal assert_dout_net_x1: std_logic_vector(8 downto 0);
  signal ce_1_sg_x119: std_logic;
  signal clk_1_sg_x119: std_logic;
  signal concat_y_net_x1: std_logic_vector(8 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x119 <= ce_1;
  clk_1_sg_x119 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_6677c7a36d: entity work.add_convert0_entity_6677c7a36d
    port map (
      ce_1 => ce_1_sg_x119,
      clk_1 => clk_1_sg_x119,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_9b7575767f: entity work.add_convert1_entity_9b7575767f
    port map (
      ce_1 => ce_1_sg_x119,
      clk_1 => clk_1_sg_x119,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 9,
      dout_width => 9
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_ef07e318f3: entity work.c_to_ri_entity_ef07e318f3
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x119,
      clk => clk_1_sg_x119,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x119,
      clk => clk_1_sg_x119,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x119,
      clk => clk_1_sg_x119,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_00bc692256: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x119,
      clk_1 => clk_1_sg_x119,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_17dc85599c: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x119,
      clk_1 => clk_1_sg_x119,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 9,
      c_width => 36,
      core_name0 => "bmg_72_e02664f04ec6e0c0",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x119,
      clk => clk_1_sg_x119,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen/ri_to_c"

entity ri_to_c_entity_5ed22bc0d3 is
  port (
    im: in std_logic_vector(17 downto 0); 
    re: in std_logic_vector(17 downto 0); 
    c: out std_logic_vector(35 downto 0)
  );
end ri_to_c_entity_5ed22bc0d3;

architecture structural of ri_to_c_entity_5ed22bc0d3 is
  signal concat_y_net_x4: std_logic_vector(35 downto 0);
  signal force_im_output_port_net: std_logic_vector(17 downto 0);
  signal force_re_output_port_net: std_logic_vector(17 downto 0);
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);

begin
  mux_y_net_x5 <= im;
  mux_y_net_x4 <= re;
  c <= concat_y_net_x4;

  concat: entity work.concat_b198bd62b0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => force_re_output_port_net,
      in1 => force_im_output_port_net,
      y => concat_y_net_x4
    );

  force_im: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x5,
      output_port => force_im_output_port_net
    );

  force_re: entity work.reinterpret_580feec131
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => mux_y_net_x4,
      output_port => force_re_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_25e5e2b7e2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_25e5e2b7e2;

architecture structural of coeff_gen_entity_25e5e2b7e2 is
  signal ce_1_sg_x120: std_logic;
  signal clk_1_sg_x120: std_logic;
  signal concat_y_net_x1: std_logic_vector(8 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(8 downto 0);

begin
  ce_1_sg_x120 <= ce_1;
  clk_1_sg_x120 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_f05b79004d: entity work.bit_reverse_entity_f05b79004d
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_8c6d36a3ce: entity work.cosin_entity_8c6d36a3ce
    port map (
      ce_1 => ce_1_sg_x120,
      clk_1 => clk_1_sg_x120,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x120,
      clk => clk_1_sg_x120,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_5ed22bc0d3: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 11,
      x_width => 12,
      y_width => 9
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct/twiddle"

entity twiddle_entity_208a25c7b7 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_208a25c7b7;

architecture structural of twiddle_entity_208a25c7b7 is
  signal ce_1_sg_x121: std_logic;
  signal clk_1_sg_x121: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x121 <= ce_1;
  clk_1_sg_x121 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_e5fd0829de: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x121,
      clk_1 => clk_1_sg_x121,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_1ff518d55f: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_bcd05ee4e4: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_56cf888bad: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_b0541e7d96: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x121,
      clk_1 => clk_1_sg_x121,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_25e5e2b7e2: entity work.coeff_gen_entity_25e5e2b7e2
    port map (
      ce_1 => ce_1_sg_x121,
      clk_1 => clk_1_sg_x121,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/butterfly_direct"

entity butterfly_direct_entity_8818464f6c is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_8818464f6c;

architecture structural of butterfly_direct_entity_8818464f6c is
  signal ce_1_sg_x122: std_logic;
  signal clk_1_sg_x122: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x122 <= ce_1;
  clk_1_sg_x122 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_277738c818: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      dout => concatenate_y_net_x3
    );

  bus_convert_43c000ec6d: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_74c9ce61ab: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_376e099b6a: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_cc02258db8: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_4c2c250372: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_5b3b5027bd: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_041fbb1680: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x122,
      clk => clk_1_sg_x122,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_0c663e3ca7: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_2a2e20cd83: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_8da134038a: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_208a25c7b7: entity work.twiddle_entity_208a25c7b7
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x122,
      clk_1 => clk_1_sg_x122,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/delay0"

entity delay0_entity_edf1e41f8f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_edf1e41f8f;

architecture structural of delay0_entity_edf1e41f8f is
  signal ce_1_sg_x123: std_logic;
  signal clk_1_sg_x123: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x123 <= ce_1;
  clk_1_sg_x123 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_faa52967c8
    port map (
      ce => ce_1_sg_x123,
      clk => clk_1_sg_x123,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_7f7cf6fbb7: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_b45e8409d5: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10/sync_delay"

entity sync_delay_entity_5655f4e8ca is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_5655f4e8ca;

architecture structural of sync_delay_entity_5655f4e8ca is
  signal ce_1_sg_x125: std_logic;
  signal clk_1_sg_x125: std_logic;
  signal constant1_op_net: std_logic_vector(3 downto 0);
  signal constant2_op_net: std_logic_vector(3 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(3 downto 0);
  signal counter_op_net: std_logic_vector(3 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x125 <= ce_1;
  clk_1_sg_x125 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_145086465d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_67ad97ca70
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_230536be32
    port map (
      ce => ce_1_sg_x125,
      clk => clk_1_sg_x125,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_4d3cfceaf4
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_d930162434
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_10"

entity fft_stage_10_entity_cbd0a7e571 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_10_entity_cbd0a7e571;

architecture structural of fft_stage_10_entity_cbd0a7e571 is
  signal ce_1_sg_x126: std_logic;
  signal clk_1_sg_x126: std_logic;
  signal counter_op_net: std_logic_vector(3 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x1: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x126 <= ce_1;
  clk_1_sg_x126 <= clk_1;
  reinterpret2_output_port_net_x0 <= in1;
  reinterpret1_output_port_net_x0 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x1 <= shift;
  delay0_q_net_x1 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x8;
  sync_out <= delay0_q_net_x2;

  butterfly_direct_8818464f6c: entity work.butterfly_direct_entity_8818464f6c
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x126,
      clk_1 => clk_1_sg_x126,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x8,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x2
    );

  counter: entity work.counter_6068817c97
    port map (
      ce => ce_1_sg_x126,
      clk => clk_1_sg_x126,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_edf1e41f8f: entity work.delay0_entity_edf1e41f8f
    port map (
      ce_1 => ce_1_sg_x126,
      clk_1 => clk_1_sg_x126,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_c86a918a84: entity work.delay0_entity_edf1e41f8f
    port map (
      ce_1 => ce_1_sg_x126,
      clk_1 => clk_1_sg_x126,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x0,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x1,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x126,
      clk => clk_1_sg_x126,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x126,
      clk => clk_1_sg_x126,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x126,
      clk => clk_1_sg_x126,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x126,
      clk => clk_1_sg_x126,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x1,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_5655f4e8ca: entity work.sync_delay_entity_5655f4e8ca
    port map (
      ce_1 => ce_1_sg_x126,
      clk_1 => clk_1_sg_x126,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_73471ba88c is
  port (
    in_x0: in std_logic_vector(9 downto 0); 
    out_x0: out std_logic_vector(9 downto 0)
  );
end bit_reverse_entity_73471ba88c;

architecture structural of bit_reverse_entity_73471ba88c is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(9 downto 0);
  signal slice_y_net_x0: std_logic_vector(9 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_e774b32dc9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_adc676fe6a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(9 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_adc676fe6a;

architecture structural of add_convert0_entity_adc676fe6a is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(9 downto 0);
  signal ce_1_sg_x153: std_logic;
  signal clk_1_sg_x153: std_logic;
  signal concat_y_net: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic_vector(9 downto 0);
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(10 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(8 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x153 <= ce_1;
  clk_1_sg_x153 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x153,
      clk => clk_1_sg_x153,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_4fd36a24a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 10,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x153,
      clk => clk_1_sg_x153,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_325391d82e
    port map (
      ce => ce_1_sg_x153,
      clk => clk_1_sg_x153,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x153,
      clk => clk_1_sg_x153,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x153,
      clk => clk_1_sg_x153,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_811dd91a3d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 11,
      y_width => 9
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 11,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 10,
      x_width => 11,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_5a11f0d343 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(9 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_5a11f0d343;

architecture structural of add_convert1_entity_5a11f0d343 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(9 downto 0);
  signal ce_1_sg_x154: std_logic;
  signal clk_1_sg_x154: std_logic;
  signal concat_y_net: std_logic_vector(10 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic_vector(9 downto 0);
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(10 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(8 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x154 <= ce_1;
  clk_1_sg_x154 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_4fd36a24a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 10,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_325391d82e
    port map (
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x154,
      clk => clk_1_sg_x154,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_811dd91a3d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 11,
      y_width => 9
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 11,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 10,
      x_width => 11,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_c1d9c53131 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(9 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_c1d9c53131;

architecture structural of cosin_entity_c1d9c53131 is
  signal assert_dout_net_x1: std_logic_vector(9 downto 0);
  signal ce_1_sg_x157: std_logic;
  signal clk_1_sg_x157: std_logic;
  signal concat_y_net_x1: std_logic_vector(9 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(9 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x157 <= ce_1;
  clk_1_sg_x157 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_adc676fe6a: entity work.add_convert0_entity_adc676fe6a
    port map (
      ce_1 => ce_1_sg_x157,
      clk_1 => clk_1_sg_x157,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_5a11f0d343: entity work.add_convert1_entity_5a11f0d343
    port map (
      ce_1 => ce_1_sg_x157,
      clk_1 => clk_1_sg_x157,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 10,
      dout_width => 10
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x157,
      clk => clk_1_sg_x157,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x157,
      clk => clk_1_sg_x157,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x157,
      clk => clk_1_sg_x157,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_0fb9b1424d: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x157,
      clk_1 => clk_1_sg_x157,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_c252936999: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x157,
      clk_1 => clk_1_sg_x157,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_astro_devel_core
    generic map (
      c_address_width_a => 10,
      c_address_width_b => 10,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_9f585cf1e3329833",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x157,
      a_clk => clk_1_sg_x157,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x157,
      b_clk => clk_1_sg_x157,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_e904669fbb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_e904669fbb;

architecture structural of coeff_gen_entity_e904669fbb is
  signal ce_1_sg_x158: std_logic;
  signal clk_1_sg_x158: std_logic;
  signal concat_y_net_x1: std_logic_vector(9 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(9 downto 0);

begin
  ce_1_sg_x158 <= ce_1;
  clk_1_sg_x158 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_73471ba88c: entity work.bit_reverse_entity_73471ba88c
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_c1d9c53131: entity work.cosin_entity_c1d9c53131
    port map (
      ce_1 => ce_1_sg_x158,
      clk_1 => clk_1_sg_x158,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x158,
      clk => clk_1_sg_x158,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_f1674bfd7d: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 11,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct/twiddle"

entity twiddle_entity_9a7a0a40d2 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_9a7a0a40d2;

architecture structural of twiddle_entity_9a7a0a40d2 is
  signal ce_1_sg_x159: std_logic;
  signal clk_1_sg_x159: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x159 <= ce_1;
  clk_1_sg_x159 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_b4330a1baf: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x159,
      clk_1 => clk_1_sg_x159,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_946cb5f2c3: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_94e68fb549: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_5b8ff89e6c: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_d439dd61e8: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x159,
      clk_1 => clk_1_sg_x159,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_e904669fbb: entity work.coeff_gen_entity_e904669fbb
    port map (
      ce_1 => ce_1_sg_x159,
      clk_1 => clk_1_sg_x159,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/butterfly_direct"

entity butterfly_direct_entity_7ecb45b533 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_7ecb45b533;

architecture structural of butterfly_direct_entity_7ecb45b533 is
  signal ce_1_sg_x160: std_logic;
  signal clk_1_sg_x160: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x160 <= ce_1;
  clk_1_sg_x160 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_1220409f89: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      dout => concatenate_y_net_x3
    );

  bus_convert_4473c75da3: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_28c648ed0b: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_b06f189437: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_22be6a3c49: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_b5286627b6: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_9b3a8fc91e: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_276721afb6: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x160,
      clk => clk_1_sg_x160,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_0fb937bb8a: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_1303120367: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_4a6e4f3003: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_9a7a0a40d2: entity work.twiddle_entity_9a7a0a40d2
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x160,
      clk_1 => clk_1_sg_x160,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/delay0"

entity delay0_entity_4fba67b40a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_4fba67b40a;

architecture structural of delay0_entity_4fba67b40a is
  signal ce_1_sg_x161: std_logic;
  signal clk_1_sg_x161: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x161 <= ce_1;
  clk_1_sg_x161 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_bdaf6c9e55
    port map (
      ce => ce_1_sg_x161,
      clk => clk_1_sg_x161,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_477e8bb284: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_68f3509dfc: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11/sync_delay"

entity sync_delay_entity_80e326ccfe is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_80e326ccfe;

architecture structural of sync_delay_entity_80e326ccfe is
  signal ce_1_sg_x163: std_logic;
  signal clk_1_sg_x163: std_logic;
  signal constant1_op_net: std_logic_vector(2 downto 0);
  signal constant2_op_net: std_logic_vector(2 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(2 downto 0);
  signal counter_op_net: std_logic_vector(2 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x163 <= ce_1;
  clk_1_sg_x163 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a1c496ea88
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_ed7367cb5c
    port map (
      ce => ce_1_sg_x163,
      clk => clk_1_sg_x163,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_8fc7f5539b
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_47b317dab6
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_11"

entity fft_stage_11_entity_baad9cfaf6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_11_entity_baad9cfaf6;

architecture structural of fft_stage_11_entity_baad9cfaf6 is
  signal ce_1_sg_x164: std_logic;
  signal clk_1_sg_x164: std_logic;
  signal counter_op_net: std_logic_vector(2 downto 0);
  signal delay0_q_net_x3: std_logic;
  signal delay0_q_net_x4: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x2: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x164 <= ce_1;
  clk_1_sg_x164 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x2 <= shift;
  delay0_q_net_x3 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x10;
  sync_out <= delay0_q_net_x4;

  butterfly_direct_7ecb45b533: entity work.butterfly_direct_entity_7ecb45b533
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x164,
      clk_1 => clk_1_sg_x164,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x10,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x4
    );

  counter: entity work.counter_191d4874ab
    port map (
      ce => ce_1_sg_x164,
      clk => clk_1_sg_x164,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_4fba67b40a: entity work.delay0_entity_4fba67b40a
    port map (
      ce_1 => ce_1_sg_x164,
      clk_1 => clk_1_sg_x164,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_388349d4b3: entity work.delay0_entity_4fba67b40a
    port map (
      ce_1 => ce_1_sg_x164,
      clk_1 => clk_1_sg_x164,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x3,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x3,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x164,
      clk => clk_1_sg_x164,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x164,
      clk => clk_1_sg_x164,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x164,
      clk => clk_1_sg_x164,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x164,
      clk => clk_1_sg_x164,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x2,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_80e326ccfe: entity work.sync_delay_entity_80e326ccfe
    port map (
      ce_1 => ce_1_sg_x164,
      clk_1 => clk_1_sg_x164,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_0ef6902281 is
  port (
    in_x0: in std_logic_vector(10 downto 0); 
    out_x0: out std_logic_vector(10 downto 0)
  );
end bit_reverse_entity_0ef6902281;

architecture structural of bit_reverse_entity_0ef6902281 is
  signal bit0_y_net: std_logic;
  signal bit10_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(10 downto 0);
  signal slice_y_net_x0: std_logic_vector(10 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit10: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit10_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_a0fa71d0d3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in10(0) => bit10_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_719717153f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(10 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_719717153f;

architecture structural of add_convert0_entity_719717153f is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal addsub_s_net: std_logic_vector(10 downto 0);
  signal assert_dout_net_x0: std_logic_vector(10 downto 0);
  signal backwards_y_net: std_logic;
  signal ce_1_sg_x191: std_logic;
  signal clk_1_sg_x191: std_logic;
  signal concat_y_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic;
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(11 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(9 downto 0);
  signal mux_y_net: std_logic_vector(10 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x191 <= ce_1;
  clk_1_sg_x191 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 11,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 10,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 12,
      core_name0 => "addsb_11_0_a2af903969f3f923",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 12,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 11
    )
    port map (
      a => constant4_op_net,
      b => new_add_y_net,
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      s => addsub5_s_net
    );

  backwards: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => backwards_y_net
    );

  concat: entity work.concat_7ad1e33701
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  constant4: entity work.constant_0604807f72
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 11,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      din => mux_y_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      d(0) => backwards_y_net,
      q(0) => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9769d05421
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  mux: entity work.mux_046d743d02
    port map (
      ce => ce_1_sg_x191,
      clk => clk_1_sg_x191,
      clr => '0',
      d0 => delay14_q_net,
      d1 => addsub_s_net,
      sel(0) => delay13_q_net,
      y => mux_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_26e4a659a1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(10 downto 0); 
    add: out std_logic_vector(9 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_26e4a659a1;

architecture structural of add_convert1_entity_26e4a659a1 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal addsub_s_net: std_logic_vector(10 downto 0);
  signal assert_dout_net_x1: std_logic_vector(10 downto 0);
  signal backwards_y_net: std_logic;
  signal ce_1_sg_x192: std_logic;
  signal clk_1_sg_x192: std_logic;
  signal concat_y_net: std_logic_vector(11 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal constant4_op_net: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal delay13_q_net: std_logic;
  signal delay14_q_net: std_logic_vector(9 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(11 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(9 downto 0);
  signal mux_y_net: std_logic_vector(10 downto 0);
  signal new_add_y_net: std_logic_vector(9 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x192 <= ce_1;
  clk_1_sg_x192 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 11,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 10,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 12,
      core_name0 => "addsb_11_0_a2af903969f3f923",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 12,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 11
    )
    port map (
      a => constant4_op_net,
      b => new_add_y_net,
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      s => addsub5_s_net
    );

  backwards: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => backwards_y_net
    );

  concat: entity work.concat_7ad1e33701
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  constant4: entity work.constant_0604807f72
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 11,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 10,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      din => mux_y_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      d(0) => backwards_y_net,
      q(0) => delay13_q_net
    );

  delay14: entity work.delay_cf4f99539f
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_9769d05421
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  mux: entity work.mux_046d743d02
    port map (
      ce => ce_1_sg_x192,
      clk => clk_1_sg_x192,
      clr => '0',
      d0 => delay14_q_net,
      d1 => addsub_s_net,
      sel(0) => delay13_q_net,
      y => mux_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 9,
      x_width => 12,
      y_width => 10
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_0db9cc5ac4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(10 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_0db9cc5ac4;

architecture structural of cosin_entity_0db9cc5ac4 is
  signal assert_dout_net_x1: std_logic_vector(10 downto 0);
  signal ce_1_sg_x195: std_logic;
  signal clk_1_sg_x195: std_logic;
  signal concat_y_net_x1: std_logic_vector(10 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(9 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(9 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x195 <= ce_1;
  clk_1_sg_x195 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_719717153f: entity work.add_convert0_entity_719717153f
    port map (
      ce_1 => ce_1_sg_x195,
      clk_1 => clk_1_sg_x195,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_26e4a659a1: entity work.add_convert1_entity_26e4a659a1
    port map (
      ce_1 => ce_1_sg_x195,
      clk_1 => clk_1_sg_x195,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 11,
      dout_width => 11
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x195,
      clk => clk_1_sg_x195,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x195,
      clk => clk_1_sg_x195,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x195,
      clk => clk_1_sg_x195,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_b4f42ae22f: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x195,
      clk_1 => clk_1_sg_x195,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_43ad1ec5fe: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x195,
      clk_1 => clk_1_sg_x195,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_astro_devel_core
    generic map (
      c_address_width_a => 10,
      c_address_width_b => 10,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_15a84ff1ccdd3419",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x195,
      a_clk => clk_1_sg_x195,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x195,
      b_clk => clk_1_sg_x195,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_29dfabea80 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_29dfabea80;

architecture structural of coeff_gen_entity_29dfabea80 is
  signal ce_1_sg_x196: std_logic;
  signal clk_1_sg_x196: std_logic;
  signal concat_y_net_x1: std_logic_vector(10 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(10 downto 0);

begin
  ce_1_sg_x196 <= ce_1;
  clk_1_sg_x196 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_0ef6902281: entity work.bit_reverse_entity_0ef6902281
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_0db9cc5ac4: entity work.cosin_entity_0db9cc5ac4
    port map (
      ce_1 => ce_1_sg_x196,
      clk_1 => clk_1_sg_x196,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x196,
      clk => clk_1_sg_x196,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_504318abcc: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 11,
      x_width => 12,
      y_width => 11
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct/twiddle"

entity twiddle_entity_17c9931b5d is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_17c9931b5d;

architecture structural of twiddle_entity_17c9931b5d is
  signal ce_1_sg_x197: std_logic;
  signal clk_1_sg_x197: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x197 <= ce_1;
  clk_1_sg_x197 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_1463e16a60: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x197,
      clk_1 => clk_1_sg_x197,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_d042645e6b: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_d3535f97ee: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_74f846cef1: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_a68aa7ed1a: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x197,
      clk_1 => clk_1_sg_x197,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_29dfabea80: entity work.coeff_gen_entity_29dfabea80
    port map (
      ce_1 => ce_1_sg_x197,
      clk_1 => clk_1_sg_x197,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/butterfly_direct"

entity butterfly_direct_entity_e0e7257227 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_e0e7257227;

architecture structural of butterfly_direct_entity_e0e7257227 is
  signal ce_1_sg_x198: std_logic;
  signal clk_1_sg_x198: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x198 <= ce_1;
  clk_1_sg_x198 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_04b892945c: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      dout => concatenate_y_net_x3
    );

  bus_convert_f3975e23d7: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_e8303a28e2: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_ad33e08c25: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_34097eecfe: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_91e3f819b9: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_07ae6229ab: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_679c36b93a: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x198,
      clk => clk_1_sg_x198,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_485f89b8f2: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_e6e656c3ba: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_1b26695bfa: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_17c9931b5d: entity work.twiddle_entity_17c9931b5d
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x198,
      clk_1 => clk_1_sg_x198,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/delay0"

entity delay0_entity_ba00f039f4 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_ba00f039f4;

architecture structural of delay0_entity_ba00f039f4 is
  signal ce_1_sg_x199: std_logic;
  signal clk_1_sg_x199: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x199 <= ce_1;
  clk_1_sg_x199 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_38898c80c0
    port map (
      ce => ce_1_sg_x199,
      clk => clk_1_sg_x199,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_09f4f858d7: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_5080d50dbc: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12/sync_delay"

entity sync_delay_entity_81ac36f52d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_81ac36f52d;

architecture structural of sync_delay_entity_81ac36f52d is
  signal ce_1_sg_x201: std_logic;
  signal clk_1_sg_x201: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x201 <= ce_1;
  clk_1_sg_x201 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_e095645f0c
    port map (
      ce => ce_1_sg_x201,
      clk => clk_1_sg_x201,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f9928864ea
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_12"

entity fft_stage_12_entity_a7c8193bef is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_12_entity_a7c8193bef;

architecture structural of fft_stage_12_entity_a7c8193bef is
  signal ce_1_sg_x202: std_logic;
  signal clk_1_sg_x202: std_logic;
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x3: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x202 <= ce_1;
  clk_1_sg_x202 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x11 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x3 <= shift;
  delay0_q_net_x5 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x8;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_e0e7257227: entity work.butterfly_direct_entity_e0e7257227
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x202,
      clk_1 => clk_1_sg_x202,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x8,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.counter_363af54ff2
    port map (
      ce => ce_1_sg_x202,
      clk => clk_1_sg_x202,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_ba00f039f4: entity work.delay0_entity_ba00f039f4
    port map (
      ce_1 => ce_1_sg_x202,
      clk_1 => clk_1_sg_x202,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_456815f62e: entity work.delay0_entity_ba00f039f4
    port map (
      ce_1 => ce_1_sg_x202,
      clk_1 => clk_1_sg_x202,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x5,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x11,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x5,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x202,
      clk => clk_1_sg_x202,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x202,
      clk => clk_1_sg_x202,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x202,
      clk => clk_1_sg_x202,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x202,
      clk => clk_1_sg_x202,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x3,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_81ac36f52d: entity work.sync_delay_entity_81ac36f52d
    port map (
      ce_1 => ce_1_sg_x202,
      clk_1 => clk_1_sg_x202,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_62a8379f4c is
  port (
    in_x0: in std_logic_vector(11 downto 0); 
    out_x0: out std_logic_vector(11 downto 0)
  );
end bit_reverse_entity_62a8379f4c;

architecture structural of bit_reverse_entity_62a8379f4c is
  signal bit0_y_net: std_logic;
  signal bit10_y_net: std_logic;
  signal bit11_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal bit8_y_net: std_logic;
  signal bit9_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(11 downto 0);
  signal slice_y_net_x0: std_logic_vector(11 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit10: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit10_y_net
    );

  bit11: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit11_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  bit8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit8_y_net
    );

  bit9: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit9_y_net
    );

  concat: entity work.concat_ef66525e56
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in10(0) => bit10_y_net,
      in11(0) => bit11_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      in8(0) => bit8_y_net,
      in9(0) => bit9_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_c257cc15eb is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(11 downto 0); 
    add: out std_logic_vector(10 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_c257cc15eb;

architecture structural of add_convert0_entity_c257cc15eb is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal addsub_s_net: std_logic_vector(11 downto 0);
  signal assert_dout_net_x0: std_logic_vector(11 downto 0);
  signal backwards_y_net: std_logic;
  signal ce_1_sg_x229: std_logic;
  signal clk_1_sg_x229: std_logic;
  signal concat_y_net: std_logic_vector(12 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal delay13_q_net: std_logic;
  signal delay14_q_net: std_logic_vector(10 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(12 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(10 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal new_add_y_net: std_logic_vector(10 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x229 <= ce_1;
  clk_1_sg_x229 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 12,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 11,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 13,
      core_name0 => "addsb_11_0_47829d325bbb998a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 13,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 12
    )
    port map (
      a => constant4_op_net,
      b => new_add_y_net,
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      s => addsub5_s_net
    );

  backwards: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => backwards_y_net
    );

  concat: entity work.concat_8503582fb5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  constant4: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 12,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 11,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      din => mux_y_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d(0) => backwards_y_net,
      q(0) => delay13_q_net
    );

  delay14: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_118109a960
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  mux: entity work.mux_efb9621913
    port map (
      ce => ce_1_sg_x229,
      clk => clk_1_sg_x229,
      clr => '0',
      d0 => delay14_q_net,
      d1 => addsub_s_net,
      sel(0) => delay13_q_net,
      y => mux_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 12,
      x_width => 13,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_7d7328b537 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(11 downto 0); 
    add: out std_logic_vector(10 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_7d7328b537;

architecture structural of add_convert1_entity_7d7328b537 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal addsub_s_net: std_logic_vector(11 downto 0);
  signal assert_dout_net_x1: std_logic_vector(11 downto 0);
  signal backwards_y_net: std_logic;
  signal ce_1_sg_x230: std_logic;
  signal clk_1_sg_x230: std_logic;
  signal concat_y_net: std_logic_vector(12 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal delay13_q_net: std_logic;
  signal delay14_q_net: std_logic_vector(10 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(12 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(10 downto 0);
  signal mux_y_net: std_logic_vector(11 downto 0);
  signal new_add_y_net: std_logic_vector(10 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x230 <= ce_1;
  clk_1_sg_x230 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub: entity work.xladdsub_fft_astro_devel_core
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 12,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 11,
      c_has_c_out => 0,
      c_latency => 1,
      c_output_width => 13,
      core_name0 => "addsb_11_0_47829d325bbb998a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 13,
      latency => 1,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 12
    )
    port map (
      a => constant4_op_net,
      b => new_add_y_net,
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      s => addsub5_s_net
    );

  backwards: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => backwards_y_net
    );

  concat: entity work.concat_8503582fb5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  constant4: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 12,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 11,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      din => mux_y_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d(0) => backwards_y_net,
      q(0) => delay13_q_net
    );

  delay14: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_118109a960
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  mux: entity work.mux_efb9621913
    port map (
      ce => ce_1_sg_x230,
      clk => clk_1_sg_x230,
      clr => '0',
      d0 => delay14_q_net,
      d1 => addsub_s_net,
      sel(0) => delay13_q_net,
      y => mux_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 13,
      y_width => 11
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 12,
      x_width => 13,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_17587054f6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(11 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_17587054f6;

architecture structural of cosin_entity_17587054f6 is
  signal assert_dout_net_x1: std_logic_vector(11 downto 0);
  signal ce_1_sg_x233: std_logic;
  signal clk_1_sg_x233: std_logic;
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant1_op_net: std_logic_vector(17 downto 0);
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(10 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(10 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x233 <= ce_1;
  clk_1_sg_x233 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_c257cc15eb: entity work.add_convert0_entity_c257cc15eb
    port map (
      ce_1 => ce_1_sg_x233,
      clk_1 => clk_1_sg_x233,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_7d7328b537: entity work.add_convert1_entity_7d7328b537
    port map (
      ce_1 => ce_1_sg_x233,
      clk_1 => clk_1_sg_x233,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 12,
      dout_width => 12
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant1: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x233,
      clk => clk_1_sg_x233,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x233,
      clk => clk_1_sg_x233,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x233,
      clk => clk_1_sg_x233,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_7ebb8ae8fd: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x233,
      clk_1 => clk_1_sg_x233,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_45ce3055b2: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x233,
      clk_1 => clk_1_sg_x233,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_fft_astro_devel_core
    generic map (
      c_address_width_a => 11,
      c_address_width_b => 11,
      c_width_a => 18,
      c_width_b => 18,
      core_name0 => "bmg_72_9d950569c0d7f9e8",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x233,
      a_clk => clk_1_sg_x233,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x233,
      b_clk => clk_1_sg_x233,
      dina => constant_op_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => constant2_op_net,
      web(0) => constant3_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_17f8dbc3dc is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_17f8dbc3dc;

architecture structural of coeff_gen_entity_17f8dbc3dc is
  signal ce_1_sg_x234: std_logic;
  signal clk_1_sg_x234: std_logic;
  signal concat_y_net_x1: std_logic_vector(11 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x234 <= ce_1;
  clk_1_sg_x234 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_62a8379f4c: entity work.bit_reverse_entity_62a8379f4c
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_17587054f6: entity work.cosin_entity_17587054f6
    port map (
      ce_1 => ce_1_sg_x234,
      clk_1 => clk_1_sg_x234,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x234,
      clk => clk_1_sg_x234,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_950db3cbf3: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 11,
      x_width => 12,
      y_width => 12
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct/twiddle"

entity twiddle_entity_7ef200185e is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_7ef200185e;

architecture structural of twiddle_entity_7ef200185e is
  signal ce_1_sg_x235: std_logic;
  signal clk_1_sg_x235: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x235 <= ce_1;
  clk_1_sg_x235 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_c18c2e1c99: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x235,
      clk_1 => clk_1_sg_x235,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_90b6ca6ae9: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_8f96bfac56: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_673c3a2414: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_6ee30b2865: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x235,
      clk_1 => clk_1_sg_x235,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_17f8dbc3dc: entity work.coeff_gen_entity_17f8dbc3dc
    port map (
      ce_1 => ce_1_sg_x235,
      clk_1 => clk_1_sg_x235,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/butterfly_direct"

entity butterfly_direct_entity_5f5fc1dc90 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_5f5fc1dc90;

architecture structural of butterfly_direct_entity_5f5fc1dc90 is
  signal ce_1_sg_x236: std_logic;
  signal clk_1_sg_x236: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x3: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x20: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x236 <= ce_1;
  clk_1_sg_x236 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x20;
  a_bw_x0 <= reinterpret2_output_port_net_x3;
  of_x0 <= reinterpret1_output_port_net_x5;
  sync_out <= delay0_q_net_x3;

  bus_add_6540ab76d4: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      dout => concatenate_y_net_x3
    );

  bus_convert_4fb58dc175: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_9d7100b1d8: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x20,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_norm0_d17a734339: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_657f226b06: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_e5d159b9ce: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x5
    );

  bus_scale_73cbc01aec: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_15e6933fd3: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x236,
      clk => clk_1_sg_x236,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x3
    );

  munge_6012ea91e5: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_448dd44078: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_fcfd4c6e74: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_7ef200185e: entity work.twiddle_entity_7ef200185e
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x236,
      clk_1 => clk_1_sg_x236,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/delay0"

entity delay0_entity_a6ee97dd99 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_a6ee97dd99;

architecture structural of delay0_entity_a6ee97dd99 is
  signal ce_1_sg_x237: std_logic;
  signal clk_1_sg_x237: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x237 <= ce_1;
  clk_1_sg_x237 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_e4b9fcaf02
    port map (
      ce => ce_1_sg_x237,
      clk => clk_1_sg_x237,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_6f86611724: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_de2e45a629: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13/sync_delay"

entity sync_delay_entity_647414f66e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_647414f66e;

architecture structural of sync_delay_entity_647414f66e is
  signal ce_1_sg_x239: std_logic;
  signal clk_1_sg_x239: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x239 <= ce_1;
  clk_1_sg_x239 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_e095645f0c
    port map (
      ce => ce_1_sg_x239,
      clk => clk_1_sg_x239,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f9928864ea
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_13"

entity fft_stage_13_entity_9b58366fb2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_13_entity_9b58366fb2;

architecture structural of fft_stage_13_entity_9b58366fb2 is
  signal ce_1_sg_x240: std_logic;
  signal clk_1_sg_x240: std_logic;
  signal counter_op_net: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x4: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x4: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x21: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x8: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x240 <= ce_1;
  clk_1_sg_x240 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x4 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x8;
  out2 <= reinterpret1_output_port_net_x21;
  sync_out <= delay0_q_net_x4;

  butterfly_direct_5f5fc1dc90: entity work.butterfly_direct_entity_5f5fc1dc90
    port map (
      a => reinterpret1_output_port_net_x6,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x240,
      clk_1 => clk_1_sg_x240,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x21,
      a_bw_x0 => reinterpret2_output_port_net_x8,
      of_x0 => reinterpret1_output_port_net_x5,
      sync_out => delay0_q_net_x4
    );

  counter: entity work.counter_223a0f3237
    port map (
      ce => ce_1_sg_x240,
      clk => clk_1_sg_x240,
      clr => '0',
      rst(0) => dsync0_q_net,
      op(0) => counter_op_net
    );

  delay0_a6ee97dd99: entity work.delay0_entity_a6ee97dd99
    port map (
      ce_1 => ce_1_sg_x240,
      clk_1 => clk_1_sg_x240,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_14c37cf076: entity work.delay0_entity_a6ee97dd99
    port map (
      ce_1 => ce_1_sg_x240,
      clk_1 => clk_1_sg_x240,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x6
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x7,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x240,
      clk => clk_1_sg_x240,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x240,
      clk => clk_1_sg_x240,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x5,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x240,
      clk => clk_1_sg_x240,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x240,
      clk => clk_1_sg_x240,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 12,
      new_msb => 12,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x4,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 1,
      y_width => 1
    )
    port map (
      x(0) => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_647414f66e: entity work.sync_delay_entity_647414f66e
    port map (
      ce_1 => ce_1_sg_x240,
      clk_1 => clk_1_sg_x240,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/butterfly_direct/twiddle/negate"

entity negate_entity_0d8c44cc35 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(17 downto 0); 
    dout: out std_logic_vector(17 downto 0)
  );
end negate_entity_0d8c44cc35;

architecture structural of negate_entity_0d8c44cc35 is
  signal ce_1_sg_x260: std_logic;
  signal clk_1_sg_x260: std_logic;
  signal neg1_op_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x260 <= ce_1;
  clk_1_sg_x260 <= clk_1;
  reinterpret2_output_port_net_x2 <= din;
  dout <= reinterpret1_output_port_net_x2;

  bussify_d29901d763: entity work.bussify_entity_7962d3f7d8
    port map (
      in1 => neg1_op_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

  debus_0dc62fb19f: entity work.a_debus_entity_7fbb8fef33
    port map (
      bus_in => reinterpret2_output_port_net_x2,
      msb_lsb_out1 => reinterpret1_output_port_net_x1
    );

  neg1: entity work.negate_155cd8ddf7
    port map (
      ce => ce_1_sg_x260,
      clk => clk_1_sg_x260,
      clr => '0',
      ip => reinterpret1_output_port_net_x1,
      op => neg1_op_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/butterfly_direct/twiddle"

entity twiddle_entity_c9edee7d91 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_c9edee7d91;

architecture structural of twiddle_entity_c9edee7d91 is
  signal ce_1_sg_x261: std_logic;
  signal clk_1_sg_x261: std_logic;
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay0_q_net_x4: std_logic_vector(35 downto 0);
  signal delay2_q_net: std_logic;
  signal delay3_q_net: std_logic_vector(17 downto 0);
  signal delay4_q_net: std_logic_vector(17 downto 0);
  signal delay5_q_net: std_logic_vector(17 downto 0);
  signal delay6_q_net: std_logic_vector(17 downto 0);
  signal delay7_q_net: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux0_y_net_x0: std_logic_vector(17 downto 0);
  signal mux1_y_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x0: std_logic;
  signal reinterpret1_output_port_net_x0: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(17 downto 0);
  signal reinterpret_out_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal slice_y_net: std_logic;

begin
  concatenate_y_net_x0 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x261 <= ce_1;
  clk_1_sg_x261 <= clk_1;
  mux_y_net_x0 <= sync_in;
  ao <= delay0_q_net_x4;
  bwo <= reinterpret_out_output_port_net_x5;
  sync_out <= delay8_q_net_x0;

  bus_create_d882c3b837: entity work.join_entity_92d8cf050f
    port map (
      in1 => mux0_y_net_x0,
      in2 => mux1_y_net_x0,
      bus_out => concatenate_y_net_x2
    );

  bus_expand_ff9ee87361: entity work.bus_expand_a_entity_b94579d477
    port map (
      bus_in => reinterpret_out_output_port_net_x1,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out2 => reinterpret2_output_port_net_x2
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      rst(0) => delay7_q_net,
      op => counter_op_net
    );

  delay0: entity work.delay_dbbe492743
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => concatenate_y_net_x0,
      q => delay0_q_net_x4
    );

  delay2: entity work.delay_43bd805056
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d(0) => slice_y_net,
      q(0) => delay2_q_net
    );

  delay3: entity work.delay_c462a80bee
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => delay6_q_net,
      q => delay3_q_net
    );

  delay4: entity work.delay_c462a80bee
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => reinterpret1_output_port_net_x2,
      q => delay4_q_net
    );

  delay5: entity work.delay_328e8ebbb5
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => reinterpret2_output_port_net_x2,
      q => delay5_q_net
    );

  delay6: entity work.delay_328e8ebbb5
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => delay6_q_net
    );

  delay7: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d(0) => mux_y_net_x0,
      q(0) => delay7_q_net
    );

  delay8: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d(0) => delay7_q_net,
      q(0) => delay8_q_net_x0
    );

  munge_in_76895dc91e: entity work.munge_a_entity_7fbc079bee
    port map (
      din => dmux0_q_net_x1,
      dout => reinterpret_out_output_port_net_x1
    );

  munge_out_71cae34c8e: entity work.munge_a_entity_7fbc079bee
    port map (
      din => concatenate_y_net_x2,
      dout => reinterpret_out_output_port_net_x5
    );

  mux0: entity work.mux_621a1c5abf
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d0 => delay5_q_net,
      d1 => delay6_q_net,
      sel(0) => slice_y_net,
      y => mux0_y_net_x0
    );

  mux1: entity work.mux_181e58d842
    port map (
      ce => ce_1_sg_x261,
      clk => clk_1_sg_x261,
      clr => '0',
      d0 => delay3_q_net,
      d1 => delay4_q_net,
      sel(0) => delay2_q_net,
      y => mux1_y_net_x0
    );

  negate_0d8c44cc35: entity work.negate_entity_0d8c44cc35
    port map (
      ce_1 => ce_1_sg_x261,
      clk_1 => clk_1_sg_x261,
      din => reinterpret2_output_port_net_x2,
      dout => reinterpret1_output_port_net_x2
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/butterfly_direct"

entity butterfly_direct_entity_9cfb41c90d is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_9cfb41c90d;

architecture structural of butterfly_direct_entity_9cfb41c90d is
  signal ce_1_sg_x262: std_logic;
  signal clk_1_sg_x262: std_logic;
  signal concat_y_net_x3: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(75 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(37 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal delay0_q_net_x4: std_logic_vector(35 downto 0);
  signal delay8_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x1: std_logic;
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal reinterpret_out_output_port_net_x5: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;

begin
  concatenate_y_net_x12 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x262 <= ce_1;
  clk_1_sg_x262 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x1 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x4;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x5;
  sync_out <= delay0_q_net_x0;

  bus_add_d3b585d91e: entity work.bus_add_entity_a60c7dc670
    port map (
      a => delay0_q_net_x4,
      b => reinterpret_out_output_port_net_x5,
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      dout => concatenate_y_net_x1
    );

  bus_convert_a2445ed3a0: entity work.bus_convert_entity_7b742cca79
    port map (
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_316148230e: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x4,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_8be0bd93b7: entity work.bus_norm0_entity_74bb60a7d0
    port map (
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_42a8bcdcf3: entity work.bus_norm1_entity_b00e4bc012
    port map (
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_2d953f9677: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x5
    );

  bus_scale_fcebb2494f: entity work.bus_scale_entity_316a2a993e
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_f44c020acc: entity work.bus_sub_entity_2680215111
    port map (
      a => delay0_q_net_x4,
      b => reinterpret_out_output_port_net_x5,
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_4822199898
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x1,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x262,
      clk => clk_1_sg_x262,
      clr => '0',
      d(0) => delay8_q_net_x0,
      q(0) => delay0_q_net_x0
    );

  munge_ad11101a42: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_28899cc845: entity work.mux_entity_e2fd897480
    port map (
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_5d96a6ca10: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_c9edee7d91: entity work.twiddle_entity_c9edee7d91
    port map (
      ai => concatenate_y_net_x12,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x262,
      clk_1 => clk_1_sg_x262,
      sync_in => mux_y_net_x1,
      ao => delay0_q_net_x4,
      bwo => reinterpret_out_output_port_net_x5,
      sync_out => delay8_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/debus_addr"

entity debus_addr_entity_4542e24fb0 is
  port (
    bus_in: in std_logic_vector(10 downto 0); 
    msb_lsb_out1: out std_logic_vector(10 downto 0)
  );
end debus_addr_entity_4542e24fb0;

architecture structural of debus_addr_entity_4542e24fb0 is
  signal reinterpret1_output_port_net_x1: std_logic_vector(10 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(10 downto 0);
  signal slice1_y_net: std_logic_vector(10 downto 0);

begin
  reinterpret1_output_port_net_x1 <= bus_in;
  msb_lsb_out1 <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_6b1adb5d55
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 10,
      x_width => 11,
      y_width => 11
    )
    port map (
      x => reinterpret1_output_port_net_x1,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/debus_din"

entity debus_din_entity_ac9caef803 is
  port (
    bus_in: in std_logic_vector(35 downto 0); 
    lsb_out1: out std_logic_vector(8 downto 0); 
    msb_out4: out std_logic_vector(8 downto 0); 
    out2: out std_logic_vector(8 downto 0); 
    out3: out std_logic_vector(8 downto 0)
  );
end debus_din_entity_ac9caef803;

architecture structural of debus_din_entity_ac9caef803 is
  signal ddin_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(8 downto 0);
  signal slice1_y_net: std_logic_vector(8 downto 0);
  signal slice2_y_net: std_logic_vector(8 downto 0);
  signal slice3_y_net: std_logic_vector(8 downto 0);
  signal slice4_y_net: std_logic_vector(8 downto 0);

begin
  ddin_q_net_x0 <= bus_in;
  lsb_out1 <= reinterpret1_output_port_net_x0;
  msb_out4 <= reinterpret4_output_port_net_x0;
  out2 <= reinterpret2_output_port_net_x0;
  out3 <= reinterpret3_output_port_net_x0;

  reinterpret1: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice2_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice3_y_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice4_y_net,
      output_port => reinterpret4_output_port_net_x0
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 8,
      x_width => 36,
      y_width => 9
    )
    port map (
      x => ddin_q_net_x0,
      y => slice1_y_net
    );

  slice2: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 17,
      x_width => 36,
      y_width => 9
    )
    port map (
      x => ddin_q_net_x0,
      y => slice2_y_net
    );

  slice3: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 26,
      x_width => 36,
      y_width => 9
    )
    port map (
      x => ddin_q_net_x0,
      y => slice3_y_net
    );

  slice4: entity work.xlslice
    generic map (
      new_lsb => 27,
      new_msb => 35,
      x_width => 36,
      y_width => 9
    )
    port map (
      x => ddin_q_net_x0,
      y => slice4_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/din_bussify"

entity din_bussify_entity_9b291bea4a is
  port (
    in1: in std_logic_vector(8 downto 0); 
    in2: in std_logic_vector(8 downto 0); 
    in3: in std_logic_vector(8 downto 0); 
    in4: in std_logic_vector(8 downto 0); 
    bus_out: out std_logic_vector(35 downto 0)
  );
end din_bussify_entity_9b291bea4a;

architecture structural of din_bussify_entity_9b291bea4a is
  signal bram0_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(8 downto 0);
  signal concatenate_y_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(8 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(8 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(8 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(8 downto 0);

begin
  bram0_data_out_net_x0 <= in1;
  bram1_data_out_net_x0 <= in2;
  bram2_data_out_net_x0 <= in3;
  bram3_data_out_net_x0 <= in4;
  bus_out <= concatenate_y_net_x0;

  concatenate: entity work.concat_88cfa744f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret1_output_port_net,
      in1 => reinterpret2_output_port_net,
      in2 => reinterpret3_output_port_net,
      in3 => reinterpret4_output_port_net,
      y => concatenate_y_net_x0
    );

  reinterpret1: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram0_data_out_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram1_data_out_net_x0,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram2_data_out_net_x0,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_b754317574
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => bram3_data_out_net_x0,
      output_port => reinterpret4_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/rep_addr/bussify"

entity bussify_entity_ea57e7ceca is
  port (
    in1: in std_logic_vector(10 downto 0); 
    bus_out: out std_logic_vector(10 downto 0)
  );
end bussify_entity_ea57e7ceca;

architecture structural of bussify_entity_ea57e7ceca is
  signal din1_0_q_net_x0: std_logic_vector(10 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(10 downto 0);

begin
  din1_0_q_net_x0 <= in1;
  bus_out <= reinterpret1_output_port_net_x2;

  reinterpret1: entity work.reinterpret_6b1adb5d55
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => din1_0_q_net_x0,
      output_port => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/rep_addr"

entity rep_addr_entity_ba3a270ee3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic_vector(10 downto 0); 
    out_x0: out std_logic_vector(10 downto 0)
  );
end rep_addr_entity_ba3a270ee3;

architecture structural of rep_addr_entity_ba3a270ee3 is
  signal addr0_op_net_x0: std_logic_vector(10 downto 0);
  signal ce_1_sg_x263: std_logic;
  signal clk_1_sg_x263: std_logic;
  signal din0_0_q_net: std_logic_vector(10 downto 0);
  signal din1_0_q_net_x0: std_logic_vector(10 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(10 downto 0);

begin
  ce_1_sg_x263 <= ce_1;
  clk_1_sg_x263 <= clk_1;
  addr0_op_net_x0 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x3;

  bussify_ea57e7ceca: entity work.bussify_entity_ea57e7ceca
    port map (
      in1 => din1_0_q_net_x0,
      bus_out => reinterpret1_output_port_net_x3
    );

  din0_0: entity work.delay_49cb1051e0
    port map (
      ce => ce_1_sg_x263,
      clk => clk_1_sg_x263,
      clr => '0',
      d => addr0_op_net_x0,
      q => din0_0_q_net
    );

  din1_0: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 11
    )
    port map (
      ce => ce_1_sg_x263,
      clk => clk_1_sg_x263,
      d => din0_0_q_net,
      en => '1',
      rst => '1',
      q => din1_0_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0/rep_we"

entity rep_we_entity_fdf8eb66bf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end rep_we_entity_fdf8eb66bf;

architecture structural of rep_we_entity_fdf8eb66bf is
  signal ce_1_sg_x264: std_logic;
  signal clk_1_sg_x264: std_logic;
  signal din0_0_q_net: std_logic;
  signal din1_0_q_net_x0: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic;
  signal we0_op_net_x0: std_logic;

begin
  ce_1_sg_x264 <= ce_1;
  clk_1_sg_x264 <= clk_1;
  we0_op_net_x0 <= in_x0;
  out_x0 <= reinterpret1_output_port_net_x2;

  bussify_4aa6ff631c: entity work.bussify_entity_ad099992fc
    port map (
      in1 => din1_0_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

  din0_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x264,
      clk => clk_1_sg_x264,
      clr => '0',
      d(0) => we0_op_net_x0,
      q(0) => din0_0_q_net
    );

  din1_0: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x264,
      clk => clk_1_sg_x264,
      clr => '0',
      d(0) => din0_0_q_net,
      q(0) => din1_0_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/delay0"

entity delay0_entity_2a3fa2bdf6 is
  port (
    addr: in std_logic_vector(10 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    we: in std_logic; 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_2a3fa2bdf6;

architecture structural of delay0_entity_2a3fa2bdf6 is
  signal addr0_op_net_x1: std_logic_vector(10 downto 0);
  signal bram0_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram1_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram2_data_out_net_x0: std_logic_vector(8 downto 0);
  signal bram3_data_out_net_x0: std_logic_vector(8 downto 0);
  signal ce_1_sg_x265: std_logic;
  signal clk_1_sg_x265: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(35 downto 0);
  signal ddin_q_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(10 downto 0);
  signal reinterpret1_output_port_net_x3: std_logic_vector(10 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic;
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(8 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(8 downto 0);
  signal slice1_y_net_x0: std_logic;
  signal we0_op_net_x1: std_logic;

begin
  addr0_op_net_x1 <= addr;
  ce_1_sg_x265 <= ce_1;
  clk_1_sg_x265 <= clk_1;
  reinterpret1_output_port_net_x8 <= din;
  we0_op_net_x1 <= we;
  dout <= concatenate_y_net_x1;

  bram0: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 11,
      c_width => 9,
      core_name0 => "bmg_72_7eed1f270da26adb",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x2,
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      data_in => reinterpret4_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram0_data_out_net_x0
    );

  bram1: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 11,
      c_width => 9,
      core_name0 => "bmg_72_7eed1f270da26adb",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x2,
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      data_in => reinterpret3_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram1_data_out_net_x0
    );

  bram2: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 11,
      c_width => 9,
      core_name0 => "bmg_72_7eed1f270da26adb",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x2,
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      data_in => reinterpret2_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram2_data_out_net_x0
    );

  bram3: entity work.xlspram_fft_astro_devel_core
    generic map (
      c_address_width => 11,
      c_width => 9,
      core_name0 => "bmg_72_7eed1f270da26adb",
      latency => 2
    )
    port map (
      addr => reinterpret1_output_port_net_x2,
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      data_in => reinterpret1_output_port_net_x0,
      en => "1",
      rst => "0",
      we(0) => slice1_y_net_x0,
      data_out => bram3_data_out_net_x0
    );

  ddin: entity work.delay_38898c80c0
    port map (
      ce => ce_1_sg_x265,
      clk => clk_1_sg_x265,
      clr => '0',
      d => reinterpret1_output_port_net_x8,
      q => ddin_q_net_x0
    );

  debus_addr_4542e24fb0: entity work.debus_addr_entity_4542e24fb0
    port map (
      bus_in => reinterpret1_output_port_net_x3,
      msb_lsb_out1 => reinterpret1_output_port_net_x2
    );

  debus_din_ac9caef803: entity work.debus_din_entity_ac9caef803
    port map (
      bus_in => ddin_q_net_x0,
      lsb_out1 => reinterpret1_output_port_net_x0,
      msb_out4 => reinterpret4_output_port_net_x0,
      out2 => reinterpret2_output_port_net_x0,
      out3 => reinterpret3_output_port_net_x0
    );

  debus_we_3bac369686: entity work.we_expand_entity_d31ff06e83
    port map (
      bus_in => reinterpret1_output_port_net_x4,
      msb_lsb_out1 => slice1_y_net_x0
    );

  din_bussify_9b291bea4a: entity work.din_bussify_entity_9b291bea4a
    port map (
      in1 => bram0_data_out_net_x0,
      in2 => bram1_data_out_net_x0,
      in3 => bram2_data_out_net_x0,
      in4 => bram3_data_out_net_x0,
      bus_out => concatenate_y_net_x1
    );

  rep_addr_ba3a270ee3: entity work.rep_addr_entity_ba3a270ee3
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      in_x0 => addr0_op_net_x1,
      out_x0 => reinterpret1_output_port_net_x3
    );

  rep_we_fdf8eb66bf: entity work.rep_we_entity_fdf8eb66bf
    port map (
      ce_1 => ce_1_sg_x265,
      clk_1 => clk_1_sg_x265,
      in_x0 => we0_op_net_x1,
      out_x0 => reinterpret1_output_port_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2/sync_delay"

entity sync_delay_entity_0f20174fac is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_0f20174fac;

architecture structural of sync_delay_entity_0f20174fac is
  signal ce_1_sg_x269: std_logic;
  signal clk_1_sg_x269: std_logic;
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(11 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x2: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x269 <= ce_1;
  clk_1_sg_x269 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x2;

  constant1: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_7c91b1b314
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_a0220fdf9f
    port map (
      ce => ce_1_sg_x269,
      clk => clk_1_sg_x269,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x2
    );

  relational: entity work.relational_d36fe12c1c
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_acb3c05dd0
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_2"

entity fft_stage_2_entity_b291c4f516 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_2_entity_b291c4f516;

architecture structural of fft_stage_2_entity_b291c4f516 is
  signal addr0_op_net_x1: std_logic_vector(10 downto 0);
  signal addr1_op_net_x1: std_logic_vector(10 downto 0);
  signal ce_1_sg_x270: std_logic;
  signal clk_1_sg_x270: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x14: std_logic_vector(35 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din1_q_net: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal dsync2_q_net: std_logic;
  signal fft_shift_net_x5: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net_x0: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x5: std_logic;
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;
  signal we0_op_net_x1: std_logic;
  signal we1_op_net_x1: std_logic;

begin
  ce_1_sg_x270 <= ce_1;
  clk_1_sg_x270 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x5 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x3;

  addr0: entity work.counter_e4b8f9ed4e
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      op => addr0_op_net_x1
    );

  addr1: entity work.counter_e4b8f9ed4e
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      op => addr1_op_net_x1
    );

  butterfly_direct_9cfb41c90d: entity work.butterfly_direct_entity_9cfb41c90d
    port map (
      a => concatenate_y_net_x14,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x270,
      clk_1 => clk_1_sg_x270,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x2,
      a_bw => reinterpret1_output_port_net_x6,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x5,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      rst(0) => dsync2_q_net,
      op => counter_op_net
    );

  delay0_2a3fa2bdf6: entity work.delay0_entity_2a3fa2bdf6
    port map (
      addr => addr0_op_net_x1,
      ce_1 => ce_1_sg_x270,
      clk_1 => clk_1_sg_x270,
      din => reinterpret1_output_port_net_x9,
      we => we0_op_net_x1,
      dout => concatenate_y_net_x1
    );

  delay1_3beaf8d022: entity work.delay0_entity_2a3fa2bdf6
    port map (
      addr => addr1_op_net_x1,
      ce_1 => ce_1_sg_x270,
      clk_1 => clk_1_sg_x270,
      din => mux1_y_net_x0,
      we => we1_op_net_x1,
      dout => concatenate_y_net_x14
    );

  din0: entity work.delay_38898c80c0
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d => reinterpret2_output_port_net_x3,
      q => din0_q_net
    );

  din1: entity work.delay_4b00a70dea
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d => din0_q_net,
      q => din1_q_net
    );

  dmux0: entity work.delay_7439478232
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dsync0: entity work.delay_e18fb31a3d
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d(0) => dsync2_q_net,
      q(0) => dsync1_q_net_x0
    );

  dsync2: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync2_q_net
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x5,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d0 => concatenate_y_net_x1,
      d1 => din1_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x270,
      clk => clk_1_sg_x270,
      clr => '0',
      d0 => din1_q_net,
      d1 => concatenate_y_net_x1,
      sel(0) => slice1_y_net,
      y => mux1_y_net_x0
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x5,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 11,
      new_msb => 11,
      x_width => 12,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_0f20174fac: entity work.sync_delay_entity_0f20174fac
    port map (
      ce_1 => ce_1_sg_x270,
      clk_1 => clk_1_sg_x270,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  we0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => we0_op_net_x1
    );

  we1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => we1_op_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_c3766db52a is
  port (
    in_x0: in std_logic_vector(1 downto 0); 
    out_x0: out std_logic_vector(1 downto 0)
  );
end bit_reverse_entity_c3766db52a;

architecture structural of bit_reverse_entity_c3766db52a is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(1 downto 0);
  signal slice_y_net_x0: std_logic_vector(1 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  concat: entity work.concat_e6f5ee726b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_94ad288a01 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(1 downto 0); 
    add: out std_logic_vector(1 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_94ad288a01;

architecture structural of add_convert0_entity_94ad288a01 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(1 downto 0);
  signal ce_1_sg_x297: std_logic;
  signal clk_1_sg_x297: std_logic;
  signal concat_y_net: std_logic_vector(2 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal delay13_q_net: std_logic_vector(1 downto 0);
  signal delay14_q_net: std_logic_vector(1 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(2 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic;
  signal new_add_y_net: std_logic_vector(1 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x297 <= ce_1;
  clk_1_sg_x297 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x297,
      clk => clk_1_sg_x297,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_6160d7387c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1(0) => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 2,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 2,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x297,
      clk => clk_1_sg_x297,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_fcebea29b9
    port map (
      ce => ce_1_sg_x297,
      clk => clk_1_sg_x297,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x297,
      clk => clk_1_sg_x297,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x297,
      clk => clk_1_sg_x297,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_4a9a9a25a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => fluff_y_net,
      y(0) => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 2,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_178db56c81 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(1 downto 0); 
    add: out std_logic_vector(1 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_178db56c81;

architecture structural of add_convert1_entity_178db56c81 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(1 downto 0);
  signal ce_1_sg_x298: std_logic;
  signal clk_1_sg_x298: std_logic;
  signal concat_y_net: std_logic_vector(2 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal delay13_q_net: std_logic_vector(1 downto 0);
  signal delay14_q_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(2 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic;
  signal new_add_y_net: std_logic_vector(1 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x298 <= ce_1;
  clk_1_sg_x298 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_6160d7387c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1(0) => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 2,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 2,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_fcebea29b9
    port map (
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ce33ca7e7
    port map (
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x298,
      clk => clk_1_sg_x298,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_4a9a9a25a3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => fluff_y_net,
      y(0) => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 2,
      x_width => 3,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_173ea049e2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(1 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_173ea049e2;

architecture structural of cosin_entity_173ea049e2 is
  signal assert_dout_net_x1: std_logic_vector(1 downto 0);
  signal ce_1_sg_x301: std_logic;
  signal clk_1_sg_x301: std_logic;
  signal concat_y_net_x1: std_logic_vector(1 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(1 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(1 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x301 <= ce_1;
  clk_1_sg_x301 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_94ad288a01: entity work.add_convert0_entity_94ad288a01
    port map (
      ce_1 => ce_1_sg_x301,
      clk_1 => clk_1_sg_x301,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_178db56c81: entity work.add_convert1_entity_178db56c81
    port map (
      ce_1 => ce_1_sg_x301,
      clk_1 => clk_1_sg_x301,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 2,
      dout_width => 2
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x301,
      clk => clk_1_sg_x301,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x301,
      clk => clk_1_sg_x301,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x301,
      clk => clk_1_sg_x301,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_ff7507eb3b: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x301,
      clk_1 => clk_1_sg_x301,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_ce021af058: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x301,
      clk_1 => clk_1_sg_x301,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_astro_devel_core
    generic map (
      addr_width => 2,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_505931c5b3ea228e",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x301,
      a_clk => clk_1_sg_x301,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x301,
      b_clk => clk_1_sg_x301,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_deb21e151d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_deb21e151d;

architecture structural of coeff_gen_entity_deb21e151d is
  signal ce_1_sg_x302: std_logic;
  signal clk_1_sg_x302: std_logic;
  signal concat_y_net_x1: std_logic_vector(1 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x302 <= ce_1;
  clk_1_sg_x302 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_c3766db52a: entity work.bit_reverse_entity_c3766db52a
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_173ea049e2: entity work.cosin_entity_173ea049e2
    port map (
      ce_1 => ce_1_sg_x302,
      clk_1 => clk_1_sg_x302,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x302,
      clk => clk_1_sg_x302,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_eb459a87dc: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 11,
      x_width => 12,
      y_width => 2
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct/twiddle"

entity twiddle_entity_893ee1b873 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_893ee1b873;

architecture structural of twiddle_entity_893ee1b873 is
  signal ce_1_sg_x303: std_logic;
  signal clk_1_sg_x303: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x303 <= ce_1;
  clk_1_sg_x303 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_80d646d9a2: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_4b78adf48e: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_2430f13781: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_c06329924e: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_351a4d3932: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_deb21e151d: entity work.coeff_gen_entity_deb21e151d
    port map (
      ce_1 => ce_1_sg_x303,
      clk_1 => clk_1_sg_x303,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/butterfly_direct"

entity butterfly_direct_entity_226f5e7d6e is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_226f5e7d6e;

architecture structural of butterfly_direct_entity_226f5e7d6e is
  signal ce_1_sg_x304: std_logic;
  signal clk_1_sg_x304: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x304 <= ce_1;
  clk_1_sg_x304 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_f7fc075054: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      dout => concatenate_y_net_x3
    );

  bus_convert_22153e48a3: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_5df5e6d22f: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_96b547d138: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_0c576702e9: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_c4765078e6: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_cf85397716: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_1cc142ab2f: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x304,
      clk => clk_1_sg_x304,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_0d6356d185: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_dc4666e352: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_f4f4dd3347: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_893ee1b873: entity work.twiddle_entity_893ee1b873
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x304,
      clk_1 => clk_1_sg_x304,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/delay0"

entity delay0_entity_57ef4e9d84 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_57ef4e9d84;

architecture structural of delay0_entity_57ef4e9d84 is
  signal ce_1_sg_x305: std_logic;
  signal clk_1_sg_x305: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x305 <= ce_1;
  clk_1_sg_x305 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_e262000247
    port map (
      ce => ce_1_sg_x305,
      clk => clk_1_sg_x305,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_ed1a9dab61: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_397e0c685c: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3/sync_delay"

entity sync_delay_entity_73e91f6762 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_73e91f6762;

architecture structural of sync_delay_entity_73e91f6762 is
  signal ce_1_sg_x307: std_logic;
  signal clk_1_sg_x307: std_logic;
  signal constant1_op_net: std_logic_vector(10 downto 0);
  signal constant2_op_net: std_logic_vector(10 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(10 downto 0);
  signal counter_op_net: std_logic_vector(10 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x307 <= ce_1;
  clk_1_sg_x307 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_a3923dd146
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_0604807f72
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_118598964d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_b5e433c475
    port map (
      ce => ce_1_sg_x307,
      clk => clk_1_sg_x307,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_2147430058
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_b4b277ae0f
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_3"

entity fft_stage_3_entity_c75cf4fea1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_3_entity_c75cf4fea1;

architecture structural of fft_stage_3_entity_c75cf4fea1 is
  signal ce_1_sg_x308: std_logic;
  signal clk_1_sg_x308: std_logic;
  signal counter_op_net: std_logic_vector(10 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x6: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic;
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x308 <= ce_1;
  clk_1_sg_x308 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x6 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x10;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_226f5e7d6e: entity work.butterfly_direct_entity_226f5e7d6e
    port map (
      a => reinterpret1_output_port_net_x8,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x308,
      clk_1 => clk_1_sg_x308,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x10,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x7,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.counter_21896c7599
    port map (
      ce => ce_1_sg_x308,
      clk => clk_1_sg_x308,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_57ef4e9d84: entity work.delay0_entity_57ef4e9d84
    port map (
      ce_1 => ce_1_sg_x308,
      clk_1 => clk_1_sg_x308,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_dc233c1259: entity work.delay0_entity_57ef4e9d84
    port map (
      ce_1 => ce_1_sg_x308,
      clk_1 => clk_1_sg_x308,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x8
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x5,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x308,
      clk => clk_1_sg_x308,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x308,
      clk => clk_1_sg_x308,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x7,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x308,
      clk => clk_1_sg_x308,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x308,
      clk => clk_1_sg_x308,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x6,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 10,
      new_msb => 10,
      x_width => 11,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_73e91f6762: entity work.sync_delay_entity_73e91f6762
    port map (
      ce_1 => ce_1_sg_x308,
      clk_1 => clk_1_sg_x308,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_5248d33105 is
  port (
    in_x0: in std_logic_vector(2 downto 0); 
    out_x0: out std_logic_vector(2 downto 0)
  );
end bit_reverse_entity_5248d33105;

architecture structural of bit_reverse_entity_5248d33105 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(2 downto 0);
  signal slice_y_net_x0: std_logic_vector(2 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 3,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  concat: entity work.concat_452c4d3410
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_48d5cc476a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(2 downto 0); 
    add: out std_logic_vector(2 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_48d5cc476a;

architecture structural of add_convert0_entity_48d5cc476a is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(2 downto 0);
  signal ce_1_sg_x335: std_logic;
  signal clk_1_sg_x335: std_logic;
  signal concat_y_net: std_logic_vector(3 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal delay13_q_net: std_logic_vector(2 downto 0);
  signal delay14_q_net: std_logic_vector(2 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(3 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(1 downto 0);
  signal new_add_y_net: std_logic_vector(2 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x335 <= ce_1;
  clk_1_sg_x335 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x335,
      clk => clk_1_sg_x335,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 3,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 3,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x335,
      clk => clk_1_sg_x335,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_6edcd04662
    port map (
      ce => ce_1_sg_x335,
      clk => clk_1_sg_x335,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x335,
      clk => clk_1_sg_x335,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x335,
      clk => clk_1_sg_x335,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_949f038a6d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 4,
      y_width => 3
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_248e36a5f1 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(2 downto 0); 
    add: out std_logic_vector(2 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_248e36a5f1;

architecture structural of add_convert1_entity_248e36a5f1 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(2 downto 0);
  signal ce_1_sg_x336: std_logic;
  signal clk_1_sg_x336: std_logic;
  signal concat_y_net: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal delay13_q_net: std_logic_vector(2 downto 0);
  signal delay14_q_net: std_logic_vector(2 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(3 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(1 downto 0);
  signal new_add_y_net: std_logic_vector(2 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x336 <= ce_1;
  clk_1_sg_x336 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_bd20dd351d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 3,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 3,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_6edcd04662
    port map (
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_54d5af2115
    port map (
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x336,
      clk => clk_1_sg_x336,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_949f038a6d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 4,
      y_width => 3
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_8f338afca8 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(2 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_8f338afca8;

architecture structural of cosin_entity_8f338afca8 is
  signal assert_dout_net_x1: std_logic_vector(2 downto 0);
  signal ce_1_sg_x339: std_logic;
  signal clk_1_sg_x339: std_logic;
  signal concat_y_net_x1: std_logic_vector(2 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(2 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(2 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x339 <= ce_1;
  clk_1_sg_x339 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_48d5cc476a: entity work.add_convert0_entity_48d5cc476a
    port map (
      ce_1 => ce_1_sg_x339,
      clk_1 => clk_1_sg_x339,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_248e36a5f1: entity work.add_convert1_entity_248e36a5f1
    port map (
      ce_1 => ce_1_sg_x339,
      clk_1 => clk_1_sg_x339,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 3,
      dout_width => 3
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x339,
      clk => clk_1_sg_x339,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x339,
      clk => clk_1_sg_x339,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x339,
      clk => clk_1_sg_x339,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_a6507900ef: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x339,
      clk_1 => clk_1_sg_x339,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_6cc4d9c242: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x339,
      clk_1 => clk_1_sg_x339,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_astro_devel_core
    generic map (
      addr_width => 3,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_d20b02a9f8239c7a",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x339,
      a_clk => clk_1_sg_x339,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x339,
      b_clk => clk_1_sg_x339,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_d12ea89fbf is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_d12ea89fbf;

architecture structural of coeff_gen_entity_d12ea89fbf is
  signal ce_1_sg_x340: std_logic;
  signal clk_1_sg_x340: std_logic;
  signal concat_y_net_x1: std_logic_vector(2 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(2 downto 0);

begin
  ce_1_sg_x340 <= ce_1;
  clk_1_sg_x340 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_5248d33105: entity work.bit_reverse_entity_5248d33105
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_8f338afca8: entity work.cosin_entity_8f338afca8
    port map (
      ce_1 => ce_1_sg_x340,
      clk_1 => clk_1_sg_x340,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x340,
      clk => clk_1_sg_x340,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_390dc972f6: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 11,
      x_width => 12,
      y_width => 3
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct/twiddle"

entity twiddle_entity_969a26889f is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_969a26889f;

architecture structural of twiddle_entity_969a26889f is
  signal ce_1_sg_x341: std_logic;
  signal clk_1_sg_x341: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x341 <= ce_1;
  clk_1_sg_x341 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_0cf374d067: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_740b441704: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_19e1b0b233: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_2bd87bb94f: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_e479d26484: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_d12ea89fbf: entity work.coeff_gen_entity_d12ea89fbf
    port map (
      ce_1 => ce_1_sg_x341,
      clk_1 => clk_1_sg_x341,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/butterfly_direct"

entity butterfly_direct_entity_bf9030fc58 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_bf9030fc58;

architecture structural of butterfly_direct_entity_bf9030fc58 is
  signal ce_1_sg_x342: std_logic;
  signal clk_1_sg_x342: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x342 <= ce_1;
  clk_1_sg_x342 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_145d434f07: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      dout => concatenate_y_net_x3
    );

  bus_convert_74e2283d55: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_e1e5a010fa: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_1f793c64d8: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_758351837e: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_c0c97c78a3: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_d4fb762921: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_cd04a7efa2: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x342,
      clk => clk_1_sg_x342,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_6eb61f997e: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_d003120c32: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_257028579d: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_969a26889f: entity work.twiddle_entity_969a26889f
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x342,
      clk_1 => clk_1_sg_x342,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/delay0"

entity delay0_entity_2f5de0b955 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_2f5de0b955;

architecture structural of delay0_entity_2f5de0b955 is
  signal ce_1_sg_x343: std_logic;
  signal clk_1_sg_x343: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x343 <= ce_1;
  clk_1_sg_x343 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_0ca3374762
    port map (
      ce => ce_1_sg_x343,
      clk => clk_1_sg_x343,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_2d9a6f3e81: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_6e9144d9d5: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4/sync_delay"

entity sync_delay_entity_8f6418833f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_8f6418833f;

architecture structural of sync_delay_entity_8f6418833f is
  signal ce_1_sg_x345: std_logic;
  signal clk_1_sg_x345: std_logic;
  signal constant1_op_net: std_logic_vector(9 downto 0);
  signal constant2_op_net: std_logic_vector(9 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(9 downto 0);
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x345 <= ce_1;
  clk_1_sg_x345 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_498bc68c14
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_fbc2f0cce1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_f1ac4bddff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_d3720c25c3
    port map (
      ce => ce_1_sg_x345,
      clk => clk_1_sg_x345,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_0ffd72e037
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_f6702ea2f7
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_4"

entity fft_stage_4_entity_383ee490b3 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_4_entity_383ee490b3;

architecture structural of fft_stage_4_entity_383ee490b3 is
  signal ce_1_sg_x346: std_logic;
  signal clk_1_sg_x346: std_logic;
  signal counter_op_net: std_logic_vector(9 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x7: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x346 <= ce_1;
  clk_1_sg_x346 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x11 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x7 <= shift;
  delay0_q_net_x6 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x8;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_bf9030fc58: entity work.butterfly_direct_entity_bf9030fc58
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x346,
      clk_1 => clk_1_sg_x346,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x8,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.counter_61242a554d
    port map (
      ce => ce_1_sg_x346,
      clk => clk_1_sg_x346,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_2f5de0b955: entity work.delay0_entity_2f5de0b955
    port map (
      ce_1 => ce_1_sg_x346,
      clk_1 => clk_1_sg_x346,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_e388047ce4: entity work.delay0_entity_2f5de0b955
    port map (
      ce_1 => ce_1_sg_x346,
      clk_1 => clk_1_sg_x346,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x7,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x11,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x6,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x346,
      clk => clk_1_sg_x346,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x346,
      clk => clk_1_sg_x346,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x346,
      clk => clk_1_sg_x346,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x346,
      clk => clk_1_sg_x346,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x7,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 9,
      new_msb => 9,
      x_width => 10,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_8f6418833f: entity work.sync_delay_entity_8f6418833f
    port map (
      ce_1 => ce_1_sg_x346,
      clk_1 => clk_1_sg_x346,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_b185c3dd1f is
  port (
    in_x0: in std_logic_vector(3 downto 0); 
    out_x0: out std_logic_vector(3 downto 0)
  );
end bit_reverse_entity_b185c3dd1f;

architecture structural of bit_reverse_entity_b185c3dd1f is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(3 downto 0);
  signal slice_y_net_x0: std_logic_vector(3 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  concat: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_1358152819 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(3 downto 0); 
    add: out std_logic_vector(3 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_1358152819;

architecture structural of add_convert0_entity_1358152819 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x373: std_logic;
  signal clk_1_sg_x373: std_logic;
  signal concat_y_net: std_logic_vector(4 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal delay13_q_net: std_logic_vector(3 downto 0);
  signal delay14_q_net: std_logic_vector(3 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(4 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(2 downto 0);
  signal new_add_y_net: std_logic_vector(3 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x373 <= ce_1;
  clk_1_sg_x373 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x373,
      clk => clk_1_sg_x373,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_8f12c32de0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 4,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 4,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x373,
      clk => clk_1_sg_x373,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_4f82bd00e5
    port map (
      ce => ce_1_sg_x373,
      clk => clk_1_sg_x373,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x373,
      clk => clk_1_sg_x373,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x373,
      clk => clk_1_sg_x373,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_cf540617d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 5,
      y_width => 3
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 5,
      y_width => 4
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 5,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_98be7cda9c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(3 downto 0); 
    add: out std_logic_vector(3 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_98be7cda9c;

architecture structural of add_convert1_entity_98be7cda9c is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(3 downto 0);
  signal ce_1_sg_x374: std_logic;
  signal clk_1_sg_x374: std_logic;
  signal concat_y_net: std_logic_vector(4 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal delay13_q_net: std_logic_vector(3 downto 0);
  signal delay14_q_net: std_logic_vector(3 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(4 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(2 downto 0);
  signal new_add_y_net: std_logic_vector(3 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x374 <= ce_1;
  clk_1_sg_x374 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_8f12c32de0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 4,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 4,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_4f82bd00e5
    port map (
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_4ca77626c8
    port map (
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x374,
      clk => clk_1_sg_x374,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_cf540617d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 5,
      y_width => 3
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 5,
      y_width => 4
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 4,
      x_width => 5,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_b54cbc9939 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(3 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_b54cbc9939;

architecture structural of cosin_entity_b54cbc9939 is
  signal assert_dout_net_x1: std_logic_vector(3 downto 0);
  signal ce_1_sg_x377: std_logic;
  signal clk_1_sg_x377: std_logic;
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(3 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(3 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x377 <= ce_1;
  clk_1_sg_x377 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_1358152819: entity work.add_convert0_entity_1358152819
    port map (
      ce_1 => ce_1_sg_x377,
      clk_1 => clk_1_sg_x377,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_98be7cda9c: entity work.add_convert1_entity_98be7cda9c
    port map (
      ce_1 => ce_1_sg_x377,
      clk_1 => clk_1_sg_x377,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 4,
      dout_width => 4
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x377,
      clk => clk_1_sg_x377,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x377,
      clk => clk_1_sg_x377,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x377,
      clk => clk_1_sg_x377,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_6c08d56c12: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x377,
      clk_1 => clk_1_sg_x377,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_31f0d4b2e2: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x377,
      clk_1 => clk_1_sg_x377,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_astro_devel_core
    generic map (
      addr_width => 4,
      c_address_width => 4,
      c_width => 18,
      core_name0 => "dmg_72_efdf1b1b05926829",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x377,
      a_clk => clk_1_sg_x377,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x377,
      b_clk => clk_1_sg_x377,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_0da504c740 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_0da504c740;

architecture structural of coeff_gen_entity_0da504c740 is
  signal ce_1_sg_x378: std_logic;
  signal clk_1_sg_x378: std_logic;
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(3 downto 0);

begin
  ce_1_sg_x378 <= ce_1;
  clk_1_sg_x378 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_b185c3dd1f: entity work.bit_reverse_entity_b185c3dd1f
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_b54cbc9939: entity work.cosin_entity_b54cbc9939
    port map (
      ce_1 => ce_1_sg_x378,
      clk_1 => clk_1_sg_x378,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x378,
      clk => clk_1_sg_x378,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_b2fa954164: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 11,
      x_width => 12,
      y_width => 4
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct/twiddle"

entity twiddle_entity_87d1fd9af9 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_87d1fd9af9;

architecture structural of twiddle_entity_87d1fd9af9 is
  signal ce_1_sg_x379: std_logic;
  signal clk_1_sg_x379: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x379 <= ce_1;
  clk_1_sg_x379 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_2d5fe9f62f: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_34d61fecd3: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_5758e7605b: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_f06d586b93: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_a6fb180443: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_0da504c740: entity work.coeff_gen_entity_0da504c740
    port map (
      ce_1 => ce_1_sg_x379,
      clk_1 => clk_1_sg_x379,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/butterfly_direct"

entity butterfly_direct_entity_59e4e269f8 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_59e4e269f8;

architecture structural of butterfly_direct_entity_59e4e269f8 is
  signal ce_1_sg_x380: std_logic;
  signal clk_1_sg_x380: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x380 <= ce_1;
  clk_1_sg_x380 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_8d078d8a82: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      dout => concatenate_y_net_x3
    );

  bus_convert_8a086f9956: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_1f4faf41b5: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_bff47f6f38: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_12e8e5744b: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_8baadb1962: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_358f154c83: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_e6dab4f0ed: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x380,
      clk => clk_1_sg_x380,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_6299da6a8f: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_7400c67c2d: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_5ece24e025: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_87d1fd9af9: entity work.twiddle_entity_87d1fd9af9
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x380,
      clk_1 => clk_1_sg_x380,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/delay0"

entity delay0_entity_e195d34d2b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_e195d34d2b;

architecture structural of delay0_entity_e195d34d2b is
  signal ce_1_sg_x381: std_logic;
  signal clk_1_sg_x381: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x381 <= ce_1;
  clk_1_sg_x381 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_1f855d073b
    port map (
      ce => ce_1_sg_x381,
      clk => clk_1_sg_x381,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_9add5edd3a: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_96d20b0c6a: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5/sync_delay"

entity sync_delay_entity_9833879a3c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_9833879a3c;

architecture structural of sync_delay_entity_9833879a3c is
  signal ce_1_sg_x383: std_logic;
  signal clk_1_sg_x383: std_logic;
  signal constant1_op_net: std_logic_vector(8 downto 0);
  signal constant2_op_net: std_logic_vector(8 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(8 downto 0);
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x383 <= ce_1;
  clk_1_sg_x383 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_fd85eb7067
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_4a391b9a0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_b4ec9de7d1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_1dea202a2f
    port map (
      ce => ce_1_sg_x383,
      clk => clk_1_sg_x383,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_6c3ee657fa
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_78eac2928d
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_5"

entity fft_stage_5_entity_3a21c034a6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_5_entity_3a21c034a6;

architecture structural of fft_stage_5_entity_3a21c034a6 is
  signal ce_1_sg_x384: std_logic;
  signal clk_1_sg_x384: std_logic;
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x8: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x384 <= ce_1;
  clk_1_sg_x384 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x8 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x10;
  sync_out <= delay0_q_net_x3;

  butterfly_direct_59e4e269f8: entity work.butterfly_direct_entity_59e4e269f8
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x384,
      clk_1 => clk_1_sg_x384,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x10,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.counter_d5d467f1b8
    port map (
      ce => ce_1_sg_x384,
      clk => clk_1_sg_x384,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_e195d34d2b: entity work.delay0_entity_e195d34d2b
    port map (
      ce_1 => ce_1_sg_x384,
      clk_1 => clk_1_sg_x384,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_d12e56d207: entity work.delay0_entity_e195d34d2b
    port map (
      ce_1 => ce_1_sg_x384,
      clk_1 => clk_1_sg_x384,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x3,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x384,
      clk => clk_1_sg_x384,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x384,
      clk => clk_1_sg_x384,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x384,
      clk => clk_1_sg_x384,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x384,
      clk => clk_1_sg_x384,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x8,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 9,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_9833879a3c: entity work.sync_delay_entity_9833879a3c
    port map (
      ce_1 => ce_1_sg_x384,
      clk_1 => clk_1_sg_x384,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_1a1bf8639e is
  port (
    in_x0: in std_logic_vector(4 downto 0); 
    out_x0: out std_logic_vector(4 downto 0)
  );
end bit_reverse_entity_1a1bf8639e;

architecture structural of bit_reverse_entity_1a1bf8639e is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(4 downto 0);
  signal slice_y_net_x0: std_logic_vector(4 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  concat: entity work.concat_2b3acb49f4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_4cb29228d0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(4 downto 0); 
    add: out std_logic_vector(4 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_4cb29228d0;

architecture structural of add_convert0_entity_4cb29228d0 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(4 downto 0);
  signal ce_1_sg_x411: std_logic;
  signal clk_1_sg_x411: std_logic;
  signal concat_y_net: std_logic_vector(5 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal delay13_q_net: std_logic_vector(4 downto 0);
  signal delay14_q_net: std_logic_vector(4 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(5 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(3 downto 0);
  signal new_add_y_net: std_logic_vector(4 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x411 <= ce_1;
  clk_1_sg_x411 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x411,
      clk => clk_1_sg_x411,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_ae3f02567e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 5,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 5,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x411,
      clk => clk_1_sg_x411,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_38f665f8aa
    port map (
      ce => ce_1_sg_x411,
      clk => clk_1_sg_x411,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x411,
      clk => clk_1_sg_x411,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x411,
      clk => clk_1_sg_x411,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_ac785d9b37
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 6,
      y_width => 4
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 6,
      y_width => 5
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 5,
      x_width => 6,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_c380bab461 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(4 downto 0); 
    add: out std_logic_vector(4 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_c380bab461;

architecture structural of add_convert1_entity_c380bab461 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(4 downto 0);
  signal ce_1_sg_x412: std_logic;
  signal clk_1_sg_x412: std_logic;
  signal concat_y_net: std_logic_vector(5 downto 0);
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal delay13_q_net: std_logic_vector(4 downto 0);
  signal delay14_q_net: std_logic_vector(4 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(5 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(3 downto 0);
  signal new_add_y_net: std_logic_vector(4 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x412 <= ce_1;
  clk_1_sg_x412 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  add <= convert2_dout_net_x0;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_ae3f02567e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 5,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 5,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay13: entity work.delay_38f665f8aa
    port map (
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_b096bcf164
    port map (
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x412,
      clk => clk_1_sg_x412,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_ac785d9b37
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 6,
      y_width => 4
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 6,
      y_width => 5
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 5,
      x_width => 6,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_603630059d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(4 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_603630059d;

architecture structural of cosin_entity_603630059d is
  signal assert_dout_net_x1: std_logic_vector(4 downto 0);
  signal ce_1_sg_x415: std_logic;
  signal clk_1_sg_x415: std_logic;
  signal concat_y_net_x1: std_logic_vector(4 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal constant2_op_net: std_logic;
  signal constant_op_net: std_logic_vector(17 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(4 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(4 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal lookup_douta_net_x0: std_logic_vector(17 downto 0);
  signal lookup_doutb_net_x0: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);

begin
  ce_1_sg_x415 <= ce_1;
  clk_1_sg_x415 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_4cb29228d0: entity work.add_convert0_entity_4cb29228d0
    port map (
      ce_1 => ce_1_sg_x415,
      clk_1 => clk_1_sg_x415,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_c380bab461: entity work.add_convert1_entity_c380bab461
    port map (
      ce_1 => ce_1_sg_x415,
      clk_1 => clk_1_sg_x415,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 5,
      dout_width => 5
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant_x0: entity work.constant_95b0f967bc
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x415,
      clk => clk_1_sg_x415,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x415,
      clk => clk_1_sg_x415,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x415,
      clk => clk_1_sg_x415,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_f0c66efd87: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x415,
      clk_1 => clk_1_sg_x415,
      in_x0 => lookup_douta_net_x0,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_e7af2230d5: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x415,
      clk_1 => clk_1_sg_x415,
      in_x0 => lookup_doutb_net_x0,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  lookup: entity work.xldpram_dist_fft_astro_devel_core
    generic map (
      addr_width => 5,
      c_address_width => 5,
      c_width => 18,
      core_name0 => "dmg_72_1c323e86177437db",
      latency => 3
    )
    port map (
      a_ce => ce_1_sg_x415,
      a_clk => clk_1_sg_x415,
      addra => convert2_dout_net_x0,
      addrb => convert2_dout_net_x1,
      b_ce => ce_1_sg_x415,
      b_clk => clk_1_sg_x415,
      dina => constant_op_net,
      ena => "1",
      enb => "1",
      wea(0) => constant2_op_net,
      douta => lookup_douta_net_x0,
      doutb => lookup_doutb_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_bcfcc2a4f0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_bcfcc2a4f0;

architecture structural of coeff_gen_entity_bcfcc2a4f0 is
  signal ce_1_sg_x416: std_logic;
  signal clk_1_sg_x416: std_logic;
  signal concat_y_net_x1: std_logic_vector(4 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(4 downto 0);

begin
  ce_1_sg_x416 <= ce_1;
  clk_1_sg_x416 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_1a1bf8639e: entity work.bit_reverse_entity_1a1bf8639e
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_603630059d: entity work.cosin_entity_603630059d
    port map (
      ce_1 => ce_1_sg_x416,
      clk_1 => clk_1_sg_x416,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x416,
      clk => clk_1_sg_x416,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_3ec0cc8d4b: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 11,
      x_width => 12,
      y_width => 5
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct/twiddle"

entity twiddle_entity_33c988aa26 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_33c988aa26;

architecture structural of twiddle_entity_33c988aa26 is
  signal ce_1_sg_x417: std_logic;
  signal clk_1_sg_x417: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x417 <= ce_1;
  clk_1_sg_x417 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_f6f061424b: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_f6b8d42bee: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_97dad5ed1d: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_0857db7488: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_fc685ea66b: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_bcfcc2a4f0: entity work.coeff_gen_entity_bcfcc2a4f0
    port map (
      ce_1 => ce_1_sg_x417,
      clk_1 => clk_1_sg_x417,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/butterfly_direct"

entity butterfly_direct_entity_c58ac97e20 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_c58ac97e20;

architecture structural of butterfly_direct_entity_c58ac97e20 is
  signal ce_1_sg_x418: std_logic;
  signal clk_1_sg_x418: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x418 <= ce_1;
  clk_1_sg_x418 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_243699b7ec: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      dout => concatenate_y_net_x3
    );

  bus_convert_872a31225a: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_b09d4c5fc4: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_4a138d2e9d: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_4daf9f8131: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_91c63db562: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_c2bd85df06: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_8245104b97: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x418,
      clk => clk_1_sg_x418,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_704a0021fa: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_277fd2a3a6: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_690d3248c2: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_33c988aa26: entity work.twiddle_entity_33c988aa26
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x418,
      clk_1 => clk_1_sg_x418,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/delay0"

entity delay0_entity_11b2b7a27c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_11b2b7a27c;

architecture structural of delay0_entity_11b2b7a27c is
  signal ce_1_sg_x419: std_logic;
  signal clk_1_sg_x419: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x419 <= ce_1;
  clk_1_sg_x419 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_c33e9b879a
    port map (
      ce => ce_1_sg_x419,
      clk => clk_1_sg_x419,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_ff592a2c9c: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_e234624651: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6/sync_delay"

entity sync_delay_entity_b0efd0ccd9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_b0efd0ccd9;

architecture structural of sync_delay_entity_b0efd0ccd9 is
  signal ce_1_sg_x421: std_logic;
  signal clk_1_sg_x421: std_logic;
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant2_op_net: std_logic_vector(7 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(7 downto 0);
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x421 <= ce_1;
  clk_1_sg_x421 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_e8aae5d3bb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_b437b02512
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_a98fb09579
    port map (
      ce => ce_1_sg_x421,
      clk => clk_1_sg_x421,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_54048c8b02
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_16235eb2bf
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_6"

entity fft_stage_6_entity_5c351c5ab0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_6_entity_5c351c5ab0;

architecture structural of fft_stage_6_entity_5c351c5ab0 is
  signal ce_1_sg_x422: std_logic;
  signal clk_1_sg_x422: std_logic;
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x9: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x422 <= ce_1;
  clk_1_sg_x422 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x11 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x9 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x8;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_c58ac97e20: entity work.butterfly_direct_entity_c58ac97e20
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x422,
      clk_1 => clk_1_sg_x422,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x8,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.counter_11ccef49a2
    port map (
      ce => ce_1_sg_x422,
      clk => clk_1_sg_x422,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_11b2b7a27c: entity work.delay0_entity_11b2b7a27c
    port map (
      ce_1 => ce_1_sg_x422,
      clk_1 => clk_1_sg_x422,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_9207690c32: entity work.delay0_entity_11b2b7a27c
    port map (
      ce_1 => ce_1_sg_x422,
      clk_1 => clk_1_sg_x422,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x5,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x11,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x422,
      clk => clk_1_sg_x422,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x422,
      clk => clk_1_sg_x422,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x422,
      clk => clk_1_sg_x422,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x422,
      clk => clk_1_sg_x422,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x9,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_b0efd0ccd9: entity work.sync_delay_entity_b0efd0ccd9
    port map (
      ce_1 => ce_1_sg_x422,
      clk_1 => clk_1_sg_x422,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_5bce5043ac is
  port (
    in_x0: in std_logic_vector(5 downto 0); 
    out_x0: out std_logic_vector(5 downto 0)
  );
end bit_reverse_entity_5bce5043ac;

architecture structural of bit_reverse_entity_5bce5043ac is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(5 downto 0);
  signal slice_y_net_x0: std_logic_vector(5 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  concat: entity work.concat_2dc093ca7a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_72f5883686 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(5 downto 0); 
    add: out std_logic_vector(5 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_72f5883686;

architecture structural of add_convert0_entity_72f5883686 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(5 downto 0);
  signal ce_1_sg_x449: std_logic;
  signal clk_1_sg_x449: std_logic;
  signal concat_y_net: std_logic_vector(6 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(5 downto 0);
  signal delay13_q_net: std_logic_vector(5 downto 0);
  signal delay14_q_net: std_logic_vector(5 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(6 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(4 downto 0);
  signal new_add_y_net: std_logic_vector(5 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x449 <= ce_1;
  clk_1_sg_x449 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x449,
      clk => clk_1_sg_x449,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_75261c7c53
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 6,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 6,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x449,
      clk => clk_1_sg_x449,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_da3bb0b159
    port map (
      ce => ce_1_sg_x449,
      clk => clk_1_sg_x449,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_0b18d34058
    port map (
      ce => ce_1_sg_x449,
      clk => clk_1_sg_x449,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x449,
      clk => clk_1_sg_x449,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 4,
      x_width => 7,
      y_width => 5
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 7,
      y_width => 6
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 7,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_eca3d94374 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(5 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_eca3d94374;

architecture structural of add_convert1_entity_eca3d94374 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(5 downto 0);
  signal ce_1_sg_x450: std_logic;
  signal clk_1_sg_x450: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(6 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x450 <= ce_1;
  clk_1_sg_x450 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x450,
      clk => clk_1_sg_x450,
      clr => '0',
      s => addsub5_s_net
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x450,
      clk => clk_1_sg_x450,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x450,
      clk => clk_1_sg_x450,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 6,
      x_width => 7,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_2e181ece19 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(5 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_2e181ece19;

architecture structural of cosin_entity_2e181ece19 is
  signal assert_dout_net_x1: std_logic_vector(5 downto 0);
  signal ce_1_sg_x453: std_logic;
  signal clk_1_sg_x453: std_logic;
  signal concat_y_net_x1: std_logic_vector(5 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(5 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x453 <= ce_1;
  clk_1_sg_x453 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_72f5883686: entity work.add_convert0_entity_72f5883686
    port map (
      ce_1 => ce_1_sg_x453,
      clk_1 => clk_1_sg_x453,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_eca3d94374: entity work.add_convert1_entity_eca3d94374
    port map (
      ce_1 => ce_1_sg_x453,
      clk_1 => clk_1_sg_x453,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 6,
      dout_width => 6
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_07bbe3060c: entity work.c_to_ri_entity_ef07e318f3
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x453,
      clk => clk_1_sg_x453,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x453,
      clk => clk_1_sg_x453,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x453,
      clk => clk_1_sg_x453,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_bef3a1284f: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x453,
      clk_1 => clk_1_sg_x453,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_e92a6eef0b: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x453,
      clk_1 => clk_1_sg_x453,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 6,
      c_width => 36,
      core_name0 => "bmg_72_5ed93725c6f3d1db",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x453,
      clk => clk_1_sg_x453,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_89bf56d91b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_89bf56d91b;

architecture structural of coeff_gen_entity_89bf56d91b is
  signal ce_1_sg_x454: std_logic;
  signal clk_1_sg_x454: std_logic;
  signal concat_y_net_x1: std_logic_vector(5 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x454 <= ce_1;
  clk_1_sg_x454 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_5bce5043ac: entity work.bit_reverse_entity_5bce5043ac
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_2e181ece19: entity work.cosin_entity_2e181ece19
    port map (
      ce_1 => ce_1_sg_x454,
      clk_1 => clk_1_sg_x454,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x454,
      clk => clk_1_sg_x454,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_61ff4ceed8: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 11,
      x_width => 12,
      y_width => 6
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct/twiddle"

entity twiddle_entity_1fa0d26c8d is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_1fa0d26c8d;

architecture structural of twiddle_entity_1fa0d26c8d is
  signal ce_1_sg_x455: std_logic;
  signal clk_1_sg_x455: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x455 <= ce_1;
  clk_1_sg_x455 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_e1324d8ad2: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_3415117149: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_8708c94cc1: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_599da765ef: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_8c050963d0: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_89bf56d91b: entity work.coeff_gen_entity_89bf56d91b
    port map (
      ce_1 => ce_1_sg_x455,
      clk_1 => clk_1_sg_x455,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/butterfly_direct"

entity butterfly_direct_entity_c0788de351 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_c0788de351;

architecture structural of butterfly_direct_entity_c0788de351 is
  signal ce_1_sg_x456: std_logic;
  signal clk_1_sg_x456: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x456 <= ce_1;
  clk_1_sg_x456 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_ac69e89bd8: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      dout => concatenate_y_net_x3
    );

  bus_convert_fff216cbbd: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_caa47cc32c: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_87f873e0fe: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_2603c508e7: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_ce94da770d: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_880003152c: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_cef7002465: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x456,
      clk => clk_1_sg_x456,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_bbca82ad5d: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_af069191b2: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_efafdf3706: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_1fa0d26c8d: entity work.twiddle_entity_1fa0d26c8d
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x456,
      clk_1 => clk_1_sg_x456,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/delay0"

entity delay0_entity_9ef26e0578 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_9ef26e0578;

architecture structural of delay0_entity_9ef26e0578 is
  signal ce_1_sg_x457: std_logic;
  signal clk_1_sg_x457: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x457 <= ce_1;
  clk_1_sg_x457 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_9b6c7a899e
    port map (
      ce => ce_1_sg_x457,
      clk => clk_1_sg_x457,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_f256843619: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_35b32cd9ac: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7/sync_delay"

entity sync_delay_entity_688af6bc8b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_688af6bc8b;

architecture structural of sync_delay_entity_688af6bc8b is
  signal ce_1_sg_x459: std_logic;
  signal clk_1_sg_x459: std_logic;
  signal constant1_op_net: std_logic_vector(6 downto 0);
  signal constant2_op_net: std_logic_vector(6 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(6 downto 0);
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x459 <= ce_1;
  clk_1_sg_x459 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_7244cd602b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_7b07120b87
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_180df391de
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_82d8714dde
    port map (
      ce => ce_1_sg_x459,
      clk => clk_1_sg_x459,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_9a3978c602
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_23065a6aa3
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_7"

entity fft_stage_7_entity_85b3711ade is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_7_entity_85b3711ade;

architecture structural of fft_stage_7_entity_85b3711ade is
  signal ce_1_sg_x460: std_logic;
  signal clk_1_sg_x460: std_logic;
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal delay0_q_net_x1: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x10: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x460 <= ce_1;
  clk_1_sg_x460 <= clk_1;
  reinterpret2_output_port_net_x7 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x10 <= shift;
  delay0_q_net_x6 <= sync;
  of_x0 <= logical1_y_net_x0;
  out1 <= reinterpret2_output_port_net_x2;
  out2 <= reinterpret1_output_port_net_x10;
  sync_out <= delay0_q_net_x1;

  butterfly_direct_c0788de351: entity work.butterfly_direct_entity_c0788de351
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x460,
      clk_1 => clk_1_sg_x460,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x10,
      a_bw_x0 => reinterpret2_output_port_net_x2,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x1
    );

  counter: entity work.counter_aaa565147f
    port map (
      ce => ce_1_sg_x460,
      clk => clk_1_sg_x460,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_9ef26e0578: entity work.delay0_entity_9ef26e0578
    port map (
      ce_1 => ce_1_sg_x460,
      clk_1 => clk_1_sg_x460,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_f308460704: entity work.delay0_entity_9ef26e0578
    port map (
      ce_1 => ce_1_sg_x460,
      clk_1 => clk_1_sg_x460,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x7,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x6,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x460,
      clk => clk_1_sg_x460,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x460,
      clk => clk_1_sg_x460,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x0
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x460,
      clk => clk_1_sg_x460,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x460,
      clk => clk_1_sg_x460,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x10,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_688af6bc8b: entity work.sync_delay_entity_688af6bc8b
    port map (
      ce_1 => ce_1_sg_x460,
      clk_1 => clk_1_sg_x460,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_9f02400e16 is
  port (
    in_x0: in std_logic_vector(6 downto 0); 
    out_x0: out std_logic_vector(6 downto 0)
  );
end bit_reverse_entity_9f02400e16;

architecture structural of bit_reverse_entity_9f02400e16 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(6 downto 0);
  signal slice_y_net_x0: std_logic_vector(6 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 7,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  concat: entity work.concat_eb5f1ca7f9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_271e7edde7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(6 downto 0); 
    add: out std_logic_vector(6 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_271e7edde7;

architecture structural of add_convert0_entity_271e7edde7 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(6 downto 0);
  signal ce_1_sg_x487: std_logic;
  signal clk_1_sg_x487: std_logic;
  signal concat_y_net: std_logic_vector(7 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(6 downto 0);
  signal delay13_q_net: std_logic_vector(6 downto 0);
  signal delay14_q_net: std_logic_vector(6 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(7 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(5 downto 0);
  signal new_add_y_net: std_logic_vector(6 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x487 <= ce_1;
  clk_1_sg_x487 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x487,
      clk => clk_1_sg_x487,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_dc245eb1d2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 7,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 7,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x487,
      clk => clk_1_sg_x487,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_8a9e828e57
    port map (
      ce => ce_1_sg_x487,
      clk => clk_1_sg_x487,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_9066adfc41
    port map (
      ce => ce_1_sg_x487,
      clk => clk_1_sg_x487,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x487,
      clk => clk_1_sg_x487,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_83e473517e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 6,
      x_width => 8,
      y_width => 7
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 7,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_ffbd609a05 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(6 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_ffbd609a05;

architecture structural of add_convert1_entity_ffbd609a05 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(6 downto 0);
  signal ce_1_sg_x488: std_logic;
  signal clk_1_sg_x488: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(7 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x488 <= ce_1;
  clk_1_sg_x488 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x488,
      clk => clk_1_sg_x488,
      clr => '0',
      s => addsub5_s_net
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x488,
      clk => clk_1_sg_x488,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x488,
      clk => clk_1_sg_x488,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_83e473517e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 7,
      x_width => 8,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_96f4d687ff is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(6 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_96f4d687ff;

architecture structural of cosin_entity_96f4d687ff is
  signal assert_dout_net_x1: std_logic_vector(6 downto 0);
  signal ce_1_sg_x491: std_logic;
  signal clk_1_sg_x491: std_logic;
  signal concat_y_net_x1: std_logic_vector(6 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(6 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x491 <= ce_1;
  clk_1_sg_x491 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_271e7edde7: entity work.add_convert0_entity_271e7edde7
    port map (
      ce_1 => ce_1_sg_x491,
      clk_1 => clk_1_sg_x491,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_ffbd609a05: entity work.add_convert1_entity_ffbd609a05
    port map (
      ce_1 => ce_1_sg_x491,
      clk_1 => clk_1_sg_x491,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 7,
      dout_width => 7
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_3380c4819d: entity work.c_to_ri_entity_ef07e318f3
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x491,
      clk => clk_1_sg_x491,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x491,
      clk => clk_1_sg_x491,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x491,
      clk => clk_1_sg_x491,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_4d514edc54: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x491,
      clk_1 => clk_1_sg_x491,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_f187b7fd13: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x491,
      clk_1 => clk_1_sg_x491,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 7,
      c_width => 36,
      core_name0 => "bmg_72_3d733db2a81768b0",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x491,
      clk => clk_1_sg_x491,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_b8680fe413 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_b8680fe413;

architecture structural of coeff_gen_entity_b8680fe413 is
  signal ce_1_sg_x492: std_logic;
  signal clk_1_sg_x492: std_logic;
  signal concat_y_net_x1: std_logic_vector(6 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(6 downto 0);

begin
  ce_1_sg_x492 <= ce_1;
  clk_1_sg_x492 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_9f02400e16: entity work.bit_reverse_entity_9f02400e16
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_96f4d687ff: entity work.cosin_entity_96f4d687ff
    port map (
      ce_1 => ce_1_sg_x492,
      clk_1 => clk_1_sg_x492,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x492,
      clk => clk_1_sg_x492,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_63cfe8319a: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 11,
      x_width => 12,
      y_width => 7
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct/twiddle"

entity twiddle_entity_ffd57ab662 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_ffd57ab662;

architecture structural of twiddle_entity_ffd57ab662 is
  signal ce_1_sg_x493: std_logic;
  signal clk_1_sg_x493: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x493 <= ce_1;
  clk_1_sg_x493 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_337d17dfa2: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_97b04f1efa: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_e600c33c27: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_bb2be20380: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_8b9d81a20a: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_b8680fe413: entity work.coeff_gen_entity_b8680fe413
    port map (
      ce_1 => ce_1_sg_x493,
      clk_1 => clk_1_sg_x493,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/butterfly_direct"

entity butterfly_direct_entity_a89390de2f is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_a89390de2f;

architecture structural of butterfly_direct_entity_a89390de2f is
  signal ce_1_sg_x494: std_logic;
  signal clk_1_sg_x494: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x0: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x494 <= ce_1;
  clk_1_sg_x494 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x1;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x0;

  bus_add_32bb760cb6: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      dout => concatenate_y_net_x3
    );

  bus_convert_c8dd2b14c0: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_2a2d1b5939: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x1
    );

  bus_norm0_bcf4ed7082: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_aee35666ec: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_58e601f504: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_a0cbf170d7: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_66f4c15e8e: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x494,
      clk => clk_1_sg_x494,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x0
    );

  munge_5feb06b256: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_a278efae0e: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_54a95a31d2: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_ffd57ab662: entity work.twiddle_entity_ffd57ab662
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x494,
      clk_1 => clk_1_sg_x494,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/delay0"

entity delay0_entity_64e8453fd7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_64e8453fd7;

architecture structural of delay0_entity_64e8453fd7 is
  signal ce_1_sg_x495: std_logic;
  signal clk_1_sg_x495: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x495 <= ce_1;
  clk_1_sg_x495 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_895e998e80
    port map (
      ce => ce_1_sg_x495,
      clk => clk_1_sg_x495,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_661a3cc8ac: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_376af11c68: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8/sync_delay"

entity sync_delay_entity_9cd27a4051 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_9cd27a4051;

architecture structural of sync_delay_entity_9cd27a4051 is
  signal ce_1_sg_x497: std_logic;
  signal clk_1_sg_x497: std_logic;
  signal constant1_op_net: std_logic_vector(5 downto 0);
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(5 downto 0);
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x497 <= ce_1;
  clk_1_sg_x497 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_7ea0f2fff7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_961b61f8a1
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_a267c870be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_9686286f74
    port map (
      ce => ce_1_sg_x497,
      clk => clk_1_sg_x497,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_931d61fb72
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_fe487ce1c7
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_8"

entity fft_stage_8_entity_b907805ce0 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_8_entity_b907805ce0;

architecture structural of fft_stage_8_entity_b907805ce0 is
  signal ce_1_sg_x498: std_logic;
  signal clk_1_sg_x498: std_logic;
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x11: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x8: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x498 <= ce_1;
  clk_1_sg_x498 <= clk_1;
  reinterpret2_output_port_net_x3 <= in1;
  reinterpret1_output_port_net_x11 <= in2;
  logical1_y_net_x1 <= of_in;
  fft_shift_net_x11 <= shift;
  delay0_q_net_x2 <= sync;
  of_x0 <= logical1_y_net_x2;
  out1 <= reinterpret2_output_port_net_x4;
  out2 <= reinterpret1_output_port_net_x8;
  sync_out <= delay0_q_net_x3;

  butterfly_direct_a89390de2f: entity work.butterfly_direct_entity_a89390de2f
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x498,
      clk_1 => clk_1_sg_x498,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x8,
      a_bw_x0 => reinterpret2_output_port_net_x4,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x3
    );

  counter: entity work.counter_7888581f80
    port map (
      ce => ce_1_sg_x498,
      clk => clk_1_sg_x498,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_64e8453fd7: entity work.delay0_entity_64e8453fd7
    port map (
      ce_1 => ce_1_sg_x498,
      clk_1 => clk_1_sg_x498,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_6ca7f1a82d: entity work.delay0_entity_64e8453fd7
    port map (
      ce_1 => ce_1_sg_x498,
      clk_1 => clk_1_sg_x498,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x3,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x11,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x2,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x498,
      clk => clk_1_sg_x498,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x498,
      clk => clk_1_sg_x498,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x498,
      clk => clk_1_sg_x498,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x498,
      clk => clk_1_sg_x498,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x11,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 6,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_9cd27a4051: entity work.sync_delay_entity_9cd27a4051
    port map (
      ce_1 => ce_1_sg_x498,
      clk_1 => clk_1_sg_x498,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/bit_reverse"

entity bit_reverse_entity_9e180f0aa1 is
  port (
    in_x0: in std_logic_vector(7 downto 0); 
    out_x0: out std_logic_vector(7 downto 0)
  );
end bit_reverse_entity_9e180f0aa1;

architecture structural of bit_reverse_entity_9e180f0aa1 is
  signal bit0_y_net: std_logic;
  signal bit1_y_net: std_logic;
  signal bit2_y_net: std_logic;
  signal bit3_y_net: std_logic;
  signal bit4_y_net: std_logic;
  signal bit5_y_net: std_logic;
  signal bit6_y_net: std_logic;
  signal bit7_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal slice_y_net_x0: std_logic_vector(7 downto 0);

begin
  slice_y_net_x0 <= in_x0;
  out_x0 <= concat_y_net_x0;

  bit0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit0_y_net
    );

  bit1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit1_y_net
    );

  bit2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit2_y_net
    );

  bit3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit3_y_net
    );

  bit4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit4_y_net
    );

  bit5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit5_y_net
    );

  bit6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit6_y_net
    );

  bit7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => slice_y_net_x0,
      y(0) => bit7_y_net
    );

  concat: entity work.concat_7673b9b993
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => bit0_y_net,
      in1(0) => bit1_y_net,
      in2(0) => bit2_y_net,
      in3(0) => bit3_y_net,
      in4(0) => bit4_y_net,
      in5(0) => bit5_y_net,
      in6(0) => bit6_y_net,
      in7(0) => bit7_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin/add_convert0"

entity add_convert0_entity_4162640b4d is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    theta: in std_logic_vector(7 downto 0); 
    add: out std_logic_vector(7 downto 0); 
    negate: out std_logic
  );
end add_convert0_entity_4162640b4d;

architecture structural of add_convert0_entity_4162640b4d is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x0: std_logic_vector(7 downto 0);
  signal ce_1_sg_x525: std_logic;
  signal clk_1_sg_x525: std_logic;
  signal concat_y_net: std_logic_vector(8 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(7 downto 0);
  signal delay13_q_net: std_logic_vector(7 downto 0);
  signal delay14_q_net: std_logic_vector(7 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(8 downto 0);
  signal invert_y_net: std_logic;
  signal lookup_y_net: std_logic_vector(6 downto 0);
  signal new_add_y_net: std_logic_vector(7 downto 0);
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x525 <= ce_1;
  clk_1_sg_x525 <= clk_1;
  assert_dout_net_x0 <= theta;
  add <= convert2_dout_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x525,
      clk => clk_1_sg_x525,
      clr => '0',
      s => addsub5_s_net
    );

  concat: entity work.concat_f62149b02a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => addsub5_s_net,
      in1 => lookup_y_net,
      y => concat_y_net
    );

  convert2: entity work.xlconvert_pipeline
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 8,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 8,
      latency => 2,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x525,
      clk => clk_1_sg_x525,
      clr => '0',
      din => delay13_q_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  delay13: entity work.delay_23f848c85b
    port map (
      ce => ce_1_sg_x525,
      clk => clk_1_sg_x525,
      clr => '0',
      d => delay14_q_net,
      q => delay13_q_net
    );

  delay14: entity work.delay_ebec135d8a
    port map (
      ce => ce_1_sg_x525,
      clk => clk_1_sg_x525,
      clr => '0',
      d => new_add_y_net,
      q => delay14_q_net
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x525,
      clk => clk_1_sg_x525,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_1ece14600f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x0,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  lookup: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 6,
      x_width => 9,
      y_width => 7
    )
    port map (
      x => fluff_y_net,
      y => lookup_y_net
    );

  new_add: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 9,
      y_width => 8
    )
    port map (
      x => concat_y_net,
      y => new_add_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 8,
      x_width => 9,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin/add_convert1"

entity add_convert1_entity_fd1aafb2c6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(7 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    negate: out std_logic
  );
end add_convert1_entity_fd1aafb2c6;

architecture structural of add_convert1_entity_fd1aafb2c6 is
  signal addsub5_s_net: std_logic_vector(1 downto 0);
  signal assert_dout_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x526: std_logic;
  signal clk_1_sg_x526: std_logic;
  signal concatenate_y_net_x1: std_logic_vector(72 downto 0);
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal direction_offset_op_net: std_logic_vector(1 downto 0);
  signal fluff_y_net: std_logic_vector(8 downto 0);
  signal invert_y_net: std_logic;
  signal pad_op_net: std_logic;
  signal quadrant_y_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x526 <= ce_1;
  clk_1_sg_x526 <= clk_1;
  concatenate_y_net_x1 <= misci;
  assert_dout_net_x1 <= theta;
  misco <= delay1_q_net_x0;
  negate <= delay2_q_net_x0;

  addsub5: entity work.addsub_5e958c86e4
    port map (
      a => direction_offset_op_net,
      b => quadrant_y_net,
      ce => ce_1_sg_x526,
      clk => clk_1_sg_x526,
      clr => '0',
      s => addsub5_s_net
    );

  delay1: entity work.delay_3ffe3e5660
    port map (
      ce => ce_1_sg_x526,
      clk => clk_1_sg_x526,
      clr => '0',
      d => concatenate_y_net_x1,
      q => delay1_q_net_x0
    );

  delay2: entity work.delay_a14e3dd1bd
    port map (
      ce => ce_1_sg_x526,
      clk => clk_1_sg_x526,
      clr => '0',
      d(0) => invert_y_net,
      q(0) => delay2_q_net_x0
    );

  direction_offset: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => direction_offset_op_net
    );

  fluff: entity work.concat_1ece14600f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => pad_op_net,
      in1 => assert_dout_net_x1,
      y => fluff_y_net
    );

  invert: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => addsub5_s_net,
      y(0) => invert_y_net
    );

  pad: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => pad_op_net
    );

  quadrant: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 8,
      x_width => 9,
      y_width => 2
    )
    port map (
      x => fluff_y_net,
      y => quadrant_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen/cosin"

entity cosin_entity_b5c9fcf404 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    theta: in std_logic_vector(7 downto 0); 
    cos: out std_logic_vector(17 downto 0); 
    misco: out std_logic_vector(72 downto 0); 
    sin: out std_logic_vector(17 downto 0)
  );
end cosin_entity_b5c9fcf404;

architecture structural of cosin_entity_b5c9fcf404 is
  signal assert_dout_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x529: std_logic;
  signal clk_1_sg_x529: std_logic;
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concatenate_y_net_x2: std_logic_vector(72 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(7 downto 0);
  signal delay10_q_net_x0: std_logic;
  signal delay1_q_net_x0: std_logic_vector(72 downto 0);
  signal delay1_q_net_x2: std_logic_vector(72 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay8_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic_vector(72 downto 0);
  signal force_im_output_port_net_x1: std_logic_vector(17 downto 0);
  signal force_re_output_port_net_x1: std_logic_vector(17 downto 0);
  signal mux_y_net_x2: std_logic_vector(17 downto 0);
  signal mux_y_net_x3: std_logic_vector(17 downto 0);
  signal rom_data_net_x0: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x529 <= ce_1;
  clk_1_sg_x529 <= clk_1;
  concatenate_y_net_x2 <= misci;
  concat_y_net_x1 <= theta;
  cos <= mux_y_net_x2;
  misco <= delay1_q_net_x2;
  sin <= mux_y_net_x3;

  add_convert0_4162640b4d: entity work.add_convert0_entity_4162640b4d
    port map (
      ce_1 => ce_1_sg_x529,
      clk_1 => clk_1_sg_x529,
      theta => assert_dout_net_x1,
      add => convert2_dout_net_x0,
      negate => delay2_q_net_x0
    );

  add_convert1_fd1aafb2c6: entity work.add_convert1_entity_fd1aafb2c6
    port map (
      ce_1 => ce_1_sg_x529,
      clk_1 => clk_1_sg_x529,
      misci => concatenate_y_net_x2,
      theta => assert_dout_net_x1,
      misco => delay1_q_net_x0,
      negate => delay2_q_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 8,
      dout_width => 8
    )
    port map (
      din => concat_y_net_x1,
      dout => assert_dout_net_x1
    );

  c_to_ri_8caf4f2528: entity work.c_to_ri_entity_ef07e318f3
    port map (
      c => rom_data_net_x0,
      im => force_im_output_port_net_x1,
      re => force_re_output_port_net_x1
    );

  delay: entity work.delay_4e7d828d94
    port map (
      ce => ce_1_sg_x529,
      clk => clk_1_sg_x529,
      clr => '0',
      d => delay1_q_net_x0,
      q => delay_q_net_x0
    );

  delay10: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x529,
      clk => clk_1_sg_x529,
      clr => '0',
      d(0) => delay2_q_net_x0,
      q(0) => delay10_q_net_x0
    );

  delay8: entity work.delay_23d71a76f2
    port map (
      ce => ce_1_sg_x529,
      clk => clk_1_sg_x529,
      clr => '0',
      d(0) => delay2_q_net_x1,
      q(0) => delay8_q_net_x0
    );

  invert0_5738b75360: entity work.invert0_entity_00bc692256
    port map (
      ce_1 => ce_1_sg_x529,
      clk_1 => clk_1_sg_x529,
      in_x0 => force_re_output_port_net_x1,
      negate_x0 => delay10_q_net_x0,
      out_x0 => mux_y_net_x2
    );

  invert1_db3186f6f9: entity work.invert1_entity_17dc85599c
    port map (
      ce_1 => ce_1_sg_x529,
      clk_1 => clk_1_sg_x529,
      in_x0 => force_im_output_port_net_x1,
      misci => delay_q_net_x0,
      negate_x0 => delay8_q_net_x0,
      misco => delay1_q_net_x2,
      out_x0 => mux_y_net_x3
    );

  rom: entity work.xlsprom_fft_astro_devel_core
    generic map (
      c_address_width => 8,
      c_width => 36,
      core_name0 => "bmg_72_618ffcc3f0781f68",
      latency => 2
    )
    port map (
      addr => convert2_dout_net_x0,
      ce => ce_1_sg_x529,
      clk => clk_1_sg_x529,
      en => "1",
      rst => "0",
      data => rom_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle/coeff_gen"

entity coeff_gen_entity_e391ec0b76 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    misci: in std_logic_vector(72 downto 0); 
    rst: in std_logic; 
    misco: out std_logic_vector(72 downto 0); 
    w: out std_logic_vector(35 downto 0)
  );
end coeff_gen_entity_e391ec0b76;

architecture structural of coeff_gen_entity_e391ec0b76 is
  signal ce_1_sg_x530: std_logic;
  signal clk_1_sg_x530: std_logic;
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal counter_op_net: std_logic_vector(11 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal mux_y_net_x1: std_logic;
  signal mux_y_net_x4: std_logic_vector(17 downto 0);
  signal mux_y_net_x5: std_logic_vector(17 downto 0);
  signal slice_y_net_x0: std_logic_vector(7 downto 0);

begin
  ce_1_sg_x530 <= ce_1;
  clk_1_sg_x530 <= clk_1;
  concatenate_y_net_x3 <= misci;
  mux_y_net_x1 <= rst;
  misco <= delay1_q_net_x3;
  w <= concat_y_net_x5;

  bit_reverse_9e180f0aa1: entity work.bit_reverse_entity_9e180f0aa1
    port map (
      in_x0 => slice_y_net_x0,
      out_x0 => concat_y_net_x1
    );

  cosin_b5c9fcf404: entity work.cosin_entity_b5c9fcf404
    port map (
      ce_1 => ce_1_sg_x530,
      clk_1 => clk_1_sg_x530,
      misci => concatenate_y_net_x3,
      theta => concat_y_net_x1,
      cos => mux_y_net_x4,
      misco => delay1_q_net_x3,
      sin => mux_y_net_x5
    );

  counter: entity work.counter_8f386731a6
    port map (
      ce => ce_1_sg_x530,
      clk => clk_1_sg_x530,
      clr => '0',
      rst(0) => mux_y_net_x1,
      op => counter_op_net
    );

  ri_to_c_cef8998723: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => mux_y_net_x5,
      re => mux_y_net_x4,
      c => concat_y_net_x5
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 11,
      x_width => 12,
      y_width => 8
    )
    port map (
      x => counter_op_net,
      y => slice_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct/twiddle"

entity twiddle_entity_a7009eb9f3 is
  port (
    ai: in std_logic_vector(35 downto 0); 
    bi: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sync_in: in std_logic; 
    ao: out std_logic_vector(35 downto 0); 
    bwo: out std_logic_vector(37 downto 0); 
    sync_out: out std_logic
  );
end twiddle_entity_a7009eb9f3;

architecture structural of twiddle_entity_a7009eb9f3 is
  signal ce_1_sg_x531: std_logic;
  signal clk_1_sg_x531: std_logic;
  signal concat_y_net_x5: std_logic_vector(35 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(72 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(37 downto 0);
  signal delay1_q_net_x3: std_logic_vector(72 downto 0);
  signal dmisc_q_net_x2: std_logic_vector(36 downto 0);
  signal dmisc_q_net_x3: std_logic_vector(36 downto 0);
  signal dmux0_q_net_x1: std_logic_vector(35 downto 0);
  signal mux_y_net_x2: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(73 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(36 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x2 <= ai;
  dmux0_q_net_x1 <= bi;
  ce_1_sg_x531 <= ce_1;
  clk_1_sg_x531 <= clk_1;
  mux_y_net_x2 <= sync_in;
  ao <= reinterpret1_output_port_net_x11;
  bwo <= concatenate_y_net_x7;
  sync_out <= slice2_y_net_x1;

  bus_convert_162e72eb1b: entity work.bus_convert_entity_e5fd0829de
    port map (
      ce_1 => ce_1_sg_x531,
      clk_1 => clk_1_sg_x531,
      din => reinterpret1_output_port_net_x10,
      misci => dmisc_q_net_x2,
      dout => concatenate_y_net_x7,
      misco => dmisc_q_net_x3
    );

  bus_create_f5773a2242: entity work.bus_create_entity_1ff518d55f
    port map (
      in1 => dmux0_q_net_x1,
      in2 => mux_y_net_x2,
      in3 => reinterpret1_output_port_net_x2,
      bus_out => concatenate_y_net_x3
    );

  bus_expand1_2431aa6240: entity work.bus_expand1_entity_bcd05ee4e4
    port map (
      bus_in => dmisc_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x11,
      msb_out2 => slice2_y_net_x1
    );

  bus_expand_7dfa66b4be: entity work.bus_expand_entity_56cf888bad
    port map (
      bus_in => delay1_q_net_x3,
      lsb_out1 => reinterpret1_output_port_net_x9,
      msb_out2 => reinterpret2_output_port_net_x3
    );

  bus_mult_c15fbcac02: entity work.bus_mult_entity_b0541e7d96
    port map (
      a => concat_y_net_x5,
      b => reinterpret2_output_port_net_x3,
      ce_1 => ce_1_sg_x531,
      clk_1 => clk_1_sg_x531,
      misci => reinterpret1_output_port_net_x9,
      a_b => reinterpret1_output_port_net_x10,
      misco => dmisc_q_net_x2
    );

  coeff_gen_e391ec0b76: entity work.coeff_gen_entity_e391ec0b76
    port map (
      ce_1 => ce_1_sg_x531,
      clk_1 => clk_1_sg_x531,
      misci => concatenate_y_net_x3,
      rst => mux_y_net_x2,
      misco => delay1_q_net_x3,
      w => concat_y_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/butterfly_direct"

entity butterfly_direct_entity_519720f7b6 is
  port (
    a: in std_logic_vector(35 downto 0); 
    b: in std_logic_vector(35 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    shift: in std_logic; 
    sync_in: in std_logic; 
    a_bw: out std_logic_vector(35 downto 0); 
    a_bw_x0: out std_logic_vector(35 downto 0); 
    of_x0: out std_logic; 
    sync_out: out std_logic
  );
end butterfly_direct_entity_519720f7b6;

architecture structural of butterfly_direct_entity_519720f7b6 is
  signal ce_1_sg_x532: std_logic;
  signal clk_1_sg_x532: std_logic;
  signal concat_y_net_x3: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x10: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x11: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x12: std_logic_vector(37 downto 0);
  signal concatenate_y_net_x3: std_logic_vector(39 downto 0);
  signal concatenate_y_net_x4: std_logic_vector(79 downto 0);
  signal concatenate_y_net_x5: std_logic_vector(71 downto 0);
  signal concatenate_y_net_x6: std_logic_vector(3 downto 0);
  signal concatenate_y_net_x7: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x8: std_logic_vector(83 downto 0);
  signal concatenate_y_net_x9: std_logic_vector(39 downto 0);
  signal constant_op_net_x1: std_logic_vector(3 downto 0);
  signal delay0_q_net_x2: std_logic;
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal mux_y_net_x3: std_logic;
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret2_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret_out_output_port_net_x2: std_logic_vector(3 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice2_y_net_x1: std_logic;

begin
  reinterpret1_output_port_net_x4 <= a;
  dmux0_q_net_x2 <= b;
  ce_1_sg_x532 <= ce_1;
  clk_1_sg_x532 <= clk_1;
  slice0_y_net_x1 <= shift;
  mux_y_net_x3 <= sync_in;
  a_bw <= reinterpret1_output_port_net_x5;
  a_bw_x0 <= reinterpret2_output_port_net_x2;
  of_x0 <= reinterpret1_output_port_net_x6;
  sync_out <= delay0_q_net_x2;

  bus_add_2933876691: entity work.bus_add_entity_277738c818
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      dout => concatenate_y_net_x3
    );

  bus_convert_3e5bd35afa: entity work.bus_convert_entity_43c000ec6d
    port map (
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      din => concatenate_y_net_x10,
      dout => concatenate_y_net_x5,
      overflow => concatenate_y_net_x6
    );

  bus_expand_49405ae0a2: entity work.bus_expand_entity_f69635d38b
    port map (
      bus_in => concatenate_y_net_x5,
      lsb_out1 => reinterpret1_output_port_net_x5,
      msb_out2 => reinterpret2_output_port_net_x2
    );

  bus_norm0_dc0c4c34ee: entity work.bus_norm0_entity_376e099b6a
    port map (
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      din => concat_y_net_x3,
      dout => concatenate_y_net_x7
    );

  bus_norm1_54841c7fd1: entity work.bus_norm1_entity_cc02258db8
    port map (
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      din => concatenate_y_net_x4,
      dout => concatenate_y_net_x8
    );

  bus_relational_f1e34b647b: entity work.bus_relational_entity_ea2675d756
    port map (
      a => constant_op_net_x1,
      b => reinterpret_out_output_port_net_x2,
      a_b => reinterpret1_output_port_net_x6
    );

  bus_scale_d2e5e37e79: entity work.bus_scale_entity_5b3b5027bd
    port map (
      din => concat_y_net_x3,
      dout => concatenate_y_net_x4
    );

  bus_sub_8bc5f8823f: entity work.bus_sub_entity_041fbb1680
    port map (
      a => reinterpret1_output_port_net_x11,
      b => concatenate_y_net_x12,
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      dout => concatenate_y_net_x9
    );

  concat: entity work.concat_cfdc93535e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concatenate_y_net_x3,
      in1 => concatenate_y_net_x9,
      y => concat_y_net_x3
    );

  constant_x0: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net_x1
    );

  delay0: entity work.delay_aab7b18c27
    port map (
      ce => ce_1_sg_x532,
      clk => clk_1_sg_x532,
      clr => '0',
      d(0) => slice2_y_net_x1,
      q(0) => delay0_q_net_x2
    );

  munge_5ab71a6b53: entity work.munge_entity_8c0725027d
    port map (
      din => concatenate_y_net_x6,
      dout => reinterpret_out_output_port_net_x2
    );

  mux_d1bfc4a63b: entity work.mux_entity_2a2e20cd83
    port map (
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      d0 => concatenate_y_net_x7,
      d1 => concatenate_y_net_x8,
      sel => concatenate_y_net_x11,
      out_x0 => concatenate_y_net_x10
    );

  shift_replicate_8e54698bab: entity work.shift_replicate_entity_a296056610
    port map (
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      in_x0 => slice0_y_net_x1,
      out_x0 => concatenate_y_net_x11
    );

  twiddle_a7009eb9f3: entity work.twiddle_entity_a7009eb9f3
    port map (
      ai => reinterpret1_output_port_net_x4,
      bi => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x532,
      clk_1 => clk_1_sg_x532,
      sync_in => mux_y_net_x3,
      ao => reinterpret1_output_port_net_x11,
      bwo => concatenate_y_net_x12,
      sync_out => slice2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/delay0"

entity delay0_entity_057bfc9f9e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(35 downto 0); 
    dout: out std_logic_vector(35 downto 0)
  );
end delay0_entity_057bfc9f9e;

architecture structural of delay0_entity_057bfc9f9e is
  signal ce_1_sg_x533: std_logic;
  signal clk_1_sg_x533: std_logic;
  signal del1_q_net_x0: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);

begin
  ce_1_sg_x533 <= ce_1;
  clk_1_sg_x533 <= clk_1;
  din2_q_net_x1 <= din;
  dout <= reinterpret1_output_port_net_x2;

  del1: entity work.delay_3a3620b5a6
    port map (
      ce => ce_1_sg_x533,
      clk => clk_1_sg_x533,
      clr => '0',
      d => reinterpret1_output_port_net_x0,
      q => del1_q_net_x0
    );

  din_expand_1e43b371ea: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => din2_q_net_x1,
      msb_lsb_out1 => reinterpret1_output_port_net_x0
    );

  dout_compress_3477fa150c: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => del1_q_net_x0,
      bus_out => reinterpret1_output_port_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9/sync_delay"

entity sync_delay_entity_f283fd0998 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in_x0: in std_logic; 
    out_x0: out std_logic
  );
end sync_delay_entity_f283fd0998;

architecture structural of sync_delay_entity_f283fd0998 is
  signal ce_1_sg_x535: std_logic;
  signal clk_1_sg_x535: std_logic;
  signal constant1_op_net: std_logic_vector(4 downto 0);
  signal constant2_op_net: std_logic_vector(4 downto 0);
  signal constant3_op_net: std_logic;
  signal constant_op_net: std_logic_vector(4 downto 0);
  signal counter_op_net: std_logic_vector(4 downto 0);
  signal dsync1_q_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net_x4: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x535 <= ce_1;
  clk_1_sg_x535 <= clk_1;
  dsync1_q_net_x0 <= in_x0;
  out_x0 <= mux_y_net_x4;

  constant1: entity work.constant_fe72737ca0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_ef0e2e5fc6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant_x0: entity work.constant_582a3706dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.counter_9e5adb68be
    port map (
      ce => ce_1_sg_x535,
      clk => clk_1_sg_x535,
      clr => '0',
      din => constant2_op_net,
      en(0) => logical_y_net,
      load(0) => dsync1_q_net_x0,
      op => counter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational1_op_net,
      y(0) => logical_y_net
    );

  mux: entity work.mux_1bef4ba0e4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => dsync1_q_net_x0,
      d1(0) => relational_op_net,
      sel(0) => constant3_op_net,
      y(0) => mux_y_net_x4
    );

  relational: entity work.relational_9ece3c8c4e
    port map (
      a => constant_op_net,
      b => counter_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_dc5bc996c9
    port map (
      a => counter_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core/fft_stage_9"

entity fft_stage_9_entity_c7e8d97b89 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    in1: in std_logic_vector(35 downto 0); 
    in2: in std_logic_vector(35 downto 0); 
    of_in: in std_logic; 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_stage_9_entity_c7e8d97b89;

architecture structural of fft_stage_9_entity_c7e8d97b89 is
  signal ce_1_sg_x536: std_logic;
  signal clk_1_sg_x536: std_logic;
  signal counter_op_net: std_logic_vector(4 downto 0);
  signal delay0_q_net_x4: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal din0_q_net: std_logic_vector(35 downto 0);
  signal din2_q_net_x1: std_logic_vector(35 downto 0);
  signal dmux0_q_net_x2: std_logic_vector(35 downto 0);
  signal dmux1_q_net_x1: std_logic_vector(35 downto 0);
  signal dsync0_q_net: std_logic;
  signal dsync1_q_net_x0: std_logic;
  signal fft_shift_net_x12: std_logic_vector(31 downto 0);
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal mux0_y_net: std_logic_vector(35 downto 0);
  signal mux1_y_net: std_logic_vector(35 downto 0);
  signal mux_y_net_x4: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x2: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic;
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal slice0_y_net_x1: std_logic;
  signal slice1_y_net: std_logic;

begin
  ce_1_sg_x536 <= ce_1;
  clk_1_sg_x536 <= clk_1;
  reinterpret2_output_port_net_x5 <= in1;
  reinterpret1_output_port_net_x9 <= in2;
  logical1_y_net_x3 <= of_in;
  fft_shift_net_x12 <= shift;
  delay0_q_net_x4 <= sync;
  of_x0 <= logical1_y_net_x4;
  out1 <= reinterpret2_output_port_net_x6;
  out2 <= reinterpret1_output_port_net_x10;
  sync_out <= delay0_q_net_x5;

  butterfly_direct_519720f7b6: entity work.butterfly_direct_entity_519720f7b6
    port map (
      a => reinterpret1_output_port_net_x7,
      b => dmux0_q_net_x2,
      ce_1 => ce_1_sg_x536,
      clk_1 => clk_1_sg_x536,
      shift => slice0_y_net_x1,
      sync_in => mux_y_net_x4,
      a_bw => reinterpret1_output_port_net_x10,
      a_bw_x0 => reinterpret2_output_port_net_x6,
      of_x0 => reinterpret1_output_port_net_x6,
      sync_out => delay0_q_net_x5
    );

  counter: entity work.counter_743b50abe9
    port map (
      ce => ce_1_sg_x536,
      clk => clk_1_sg_x536,
      clr => '0',
      rst(0) => dsync0_q_net,
      op => counter_op_net
    );

  delay0_057bfc9f9e: entity work.delay0_entity_057bfc9f9e
    port map (
      ce_1 => ce_1_sg_x536,
      clk_1 => clk_1_sg_x536,
      din => din2_q_net_x1,
      dout => reinterpret1_output_port_net_x2
    );

  delay1_f6888c7abd: entity work.delay0_entity_057bfc9f9e
    port map (
      ce_1 => ce_1_sg_x536,
      clk_1 => clk_1_sg_x536,
      din => dmux1_q_net_x1,
      dout => reinterpret1_output_port_net_x7
    );

  din0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret2_output_port_net_x5,
      q => din0_q_net
    );

  din2: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => reinterpret1_output_port_net_x9,
      q => din2_q_net_x1
    );

  dmux0: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux0_y_net,
      q => dmux0_q_net_x2
    );

  dmux1: entity work.delay_0c0a0420a6
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => mux1_y_net,
      q => dmux1_q_net_x1
    );

  dsync0: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay0_q_net_x4,
      q(0) => dsync0_q_net
    );

  dsync1: entity work.delay_9f02caa990
    port map (
      ce => ce_1_sg_x536,
      clk => clk_1_sg_x536,
      clr => '0',
      d(0) => dsync0_q_net,
      q(0) => dsync1_q_net_x0
    );

  logical1: entity work.logical_0309b30f97
    port map (
      ce => ce_1_sg_x536,
      clk => clk_1_sg_x536,
      clr => '0',
      d0(0) => reinterpret1_output_port_net_x6,
      d1(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x4
    );

  mux0: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x536,
      clk => clk_1_sg_x536,
      clr => '0',
      d0 => reinterpret1_output_port_net_x2,
      d1 => din0_q_net,
      sel(0) => slice1_y_net,
      y => mux0_y_net
    );

  mux1: entity work.mux_4bb6f691f7
    port map (
      ce => ce_1_sg_x536,
      clk => clk_1_sg_x536,
      clr => '0',
      d0 => din0_q_net,
      d1 => reinterpret1_output_port_net_x2,
      sel(0) => slice1_y_net,
      y => mux1_y_net
    );

  slice0: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 8,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => fft_shift_net_x12,
      y(0) => slice0_y_net_x1
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 5,
      y_width => 1
    )
    port map (
      x => counter_op_net,
      y(0) => slice1_y_net
    );

  sync_delay_f283fd0998: entity work.sync_delay_entity_f283fd0998
    port map (
      ce_1 => ce_1_sg_x536,
      clk_1 => clk_1_sg_x536,
      in_x0 => dsync1_q_net_x0,
      out_x0 => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x/biplex_core"

entity biplex_core_entity_07162b7c67 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    pol1: in std_logic_vector(35 downto 0); 
    pol2: in std_logic_vector(35 downto 0); 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    out1: out std_logic_vector(35 downto 0); 
    out2: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end biplex_core_entity_07162b7c67;

architecture structural of biplex_core_entity_07162b7c67 is
  signal ce_1_sg_x537: std_logic;
  signal clk_1_sg_x537: std_logic;
  signal constant_op_net_x0: std_logic;
  signal delay0_q_net_x10: std_logic;
  signal delay0_q_net_x11: std_logic;
  signal delay0_q_net_x12: std_logic;
  signal delay0_q_net_x13: std_logic;
  signal delay0_q_net_x14: std_logic;
  signal delay0_q_net_x15: std_logic;
  signal delay0_q_net_x2: std_logic;
  signal delay0_q_net_x3: std_logic;
  signal delay0_q_net_x5: std_logic;
  signal delay0_q_net_x6: std_logic;
  signal delay0_q_net_x7: std_logic;
  signal delay0_q_net_x8: std_logic;
  signal delay0_q_net_x9: std_logic;
  signal fft_shift_net_x13: std_logic_vector(31 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x10: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x12: std_logic;
  signal logical1_y_net_x13: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical1_y_net_x7: std_logic;
  signal logical1_y_net_x8: std_logic;
  signal logical1_y_net_x9: std_logic;
  signal reinterpret1_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x13: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x17: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x18: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x19: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x22: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x23: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x24: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x25: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x9: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x10: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x11: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x12: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x13: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x14: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x15: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x16: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x9: std_logic_vector(35 downto 0);
  signal sync_net_x1: std_logic;

begin
  ce_1_sg_x537 <= ce_1;
  clk_1_sg_x537 <= clk_1;
  reinterpret1_output_port_net_x23 <= pol1;
  reinterpret1_output_port_net_x24 <= pol2;
  fft_shift_net_x13 <= shift;
  sync_net_x1 <= sync;
  of_x0 <= logical1_y_net_x13;
  out1 <= reinterpret2_output_port_net_x16;
  out2 <= reinterpret1_output_port_net_x25;
  sync_out <= delay0_q_net_x15;

  constant_x0: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net_x0
    );

  fft_stage_10_cbd0a7e571: entity work.fft_stage_10_entity_cbd0a7e571
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x6,
      in2 => reinterpret1_output_port_net_x22,
      of_in => logical1_y_net_x12,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x14,
      of_x0 => logical1_y_net_x3,
      out1 => reinterpret2_output_port_net_x4,
      out2 => reinterpret1_output_port_net_x10,
      sync_out => delay0_q_net_x3
    );

  fft_stage_11_baad9cfaf6: entity work.fft_stage_11_entity_baad9cfaf6
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x4,
      in2 => reinterpret1_output_port_net_x10,
      of_in => logical1_y_net_x3,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x3,
      of_x0 => logical1_y_net_x2,
      out1 => reinterpret2_output_port_net_x5,
      out2 => reinterpret1_output_port_net_x11,
      sync_out => delay0_q_net_x5
    );

  fft_stage_12_a7c8193bef: entity work.fft_stage_12_entity_a7c8193bef
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x5,
      in2 => reinterpret1_output_port_net_x11,
      of_in => logical1_y_net_x2,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x5,
      of_x0 => logical1_y_net_x4,
      out1 => reinterpret2_output_port_net_x7,
      out2 => reinterpret1_output_port_net_x12,
      sync_out => delay0_q_net_x6
    );

  fft_stage_13_9b58366fb2: entity work.fft_stage_13_entity_9b58366fb2
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x7,
      in2 => reinterpret1_output_port_net_x12,
      of_in => logical1_y_net_x4,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x6,
      of_x0 => logical1_y_net_x13,
      out1 => reinterpret2_output_port_net_x16,
      out2 => reinterpret1_output_port_net_x25,
      sync_out => delay0_q_net_x15
    );

  fft_stage_1_f280a22ded: entity work.fft_stage_1_entity_f280a22ded
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret1_output_port_net_x23,
      in2 => reinterpret1_output_port_net_x24,
      of_in => constant_op_net_x0,
      shift => fft_shift_net_x13,
      sync => sync_net_x1,
      of_x0 => logical1_y_net_x1,
      out1 => reinterpret2_output_port_net_x3,
      out2 => reinterpret1_output_port_net_x9,
      sync_out => delay0_q_net_x2
    );

  fft_stage_2_b291c4f516: entity work.fft_stage_2_entity_b291c4f516
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x3,
      in2 => reinterpret1_output_port_net_x9,
      of_in => logical1_y_net_x1,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x2,
      of_x0 => logical1_y_net_x5,
      out1 => reinterpret2_output_port_net_x9,
      out2 => reinterpret1_output_port_net_x13,
      sync_out => delay0_q_net_x7
    );

  fft_stage_3_c75cf4fea1: entity work.fft_stage_3_entity_c75cf4fea1
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x9,
      in2 => reinterpret1_output_port_net_x13,
      of_in => logical1_y_net_x5,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x7,
      of_x0 => logical1_y_net_x6,
      out1 => reinterpret2_output_port_net_x10,
      out2 => reinterpret1_output_port_net_x14,
      sync_out => delay0_q_net_x8
    );

  fft_stage_4_383ee490b3: entity work.fft_stage_4_entity_383ee490b3
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x10,
      in2 => reinterpret1_output_port_net_x14,
      of_in => logical1_y_net_x6,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x8,
      of_x0 => logical1_y_net_x7,
      out1 => reinterpret2_output_port_net_x11,
      out2 => reinterpret1_output_port_net_x15,
      sync_out => delay0_q_net_x9
    );

  fft_stage_5_3a21c034a6: entity work.fft_stage_5_entity_3a21c034a6
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x11,
      in2 => reinterpret1_output_port_net_x15,
      of_in => logical1_y_net_x7,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x9,
      of_x0 => logical1_y_net_x8,
      out1 => reinterpret2_output_port_net_x12,
      out2 => reinterpret1_output_port_net_x16,
      sync_out => delay0_q_net_x10
    );

  fft_stage_6_5c351c5ab0: entity work.fft_stage_6_entity_5c351c5ab0
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x12,
      in2 => reinterpret1_output_port_net_x16,
      of_in => logical1_y_net_x8,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x10,
      of_x0 => logical1_y_net_x9,
      out1 => reinterpret2_output_port_net_x13,
      out2 => reinterpret1_output_port_net_x17,
      sync_out => delay0_q_net_x11
    );

  fft_stage_7_85b3711ade: entity work.fft_stage_7_entity_85b3711ade
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x13,
      in2 => reinterpret1_output_port_net_x17,
      of_in => logical1_y_net_x9,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x11,
      of_x0 => logical1_y_net_x10,
      out1 => reinterpret2_output_port_net_x14,
      out2 => reinterpret1_output_port_net_x18,
      sync_out => delay0_q_net_x12
    );

  fft_stage_8_b907805ce0: entity work.fft_stage_8_entity_b907805ce0
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x14,
      in2 => reinterpret1_output_port_net_x18,
      of_in => logical1_y_net_x10,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x12,
      of_x0 => logical1_y_net_x11,
      out1 => reinterpret2_output_port_net_x15,
      out2 => reinterpret1_output_port_net_x19,
      sync_out => delay0_q_net_x13
    );

  fft_stage_9_c7e8d97b89: entity work.fft_stage_9_entity_c7e8d97b89
    port map (
      ce_1 => ce_1_sg_x537,
      clk_1 => clk_1_sg_x537,
      in1 => reinterpret2_output_port_net_x15,
      in2 => reinterpret1_output_port_net_x19,
      of_in => logical1_y_net_x11,
      shift => fft_shift_net_x13,
      sync => delay0_q_net_x13,
      of_x0 => logical1_y_net_x12,
      out1 => reinterpret2_output_port_net_x6,
      out2 => reinterpret1_output_port_net_x22,
      sync_out => delay0_q_net_x14
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core/fft_biplex_real_4x"

entity fft_biplex_real_4x_entity_f257ec0d37 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    pol0_in: in std_logic_vector(17 downto 0); 
    pol1_in: in std_logic_vector(17 downto 0); 
    pol2_in: in std_logic_vector(17 downto 0); 
    pol3_in: in std_logic_vector(17 downto 0); 
    shift: in std_logic_vector(31 downto 0); 
    sync: in std_logic; 
    of_x0: out std_logic; 
    pol0_out: out std_logic_vector(35 downto 0); 
    pol1_out: out std_logic_vector(35 downto 0); 
    pol2_out: out std_logic_vector(35 downto 0); 
    pol3_out: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_biplex_real_4x_entity_f257ec0d37;

architecture structural of fft_biplex_real_4x_entity_f257ec0d37 is
  signal ce_1_sg_x538: std_logic;
  signal clk_1_sg_x538: std_logic;
  signal concat_y_net_x1: std_logic_vector(35 downto 0);
  signal concat_y_net_x2: std_logic_vector(35 downto 0);
  signal delay0_q_net_x15: std_logic;
  signal fft_shift_net_x14: std_logic_vector(31 downto 0);
  signal logical1_y_net_x14: std_logic;
  signal pol1_net_x1: std_logic_vector(17 downto 0);
  signal pol2_net_x1: std_logic_vector(17 downto 0);
  signal pol3_net_x1: std_logic_vector(17 downto 0);
  signal pol4_net_x1: std_logic_vector(17 downto 0);
  signal reinterpret1_output_port_net_x20: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x21: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x22: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x23: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x24: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x25: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x26: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x4: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x5: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x6: std_logic_vector(35 downto 0);
  signal reinterpret1_output_port_net_x7: std_logic_vector(35 downto 0);
  signal reinterpret2_output_port_net_x16: std_logic_vector(35 downto 0);
  signal sync_delay1_q_net_x2: std_logic;
  signal sync_net_x2: std_logic;

begin
  ce_1_sg_x538 <= ce_1;
  clk_1_sg_x538 <= clk_1;
  pol1_net_x1 <= pol0_in;
  pol2_net_x1 <= pol1_in;
  pol3_net_x1 <= pol2_in;
  pol4_net_x1 <= pol3_in;
  fft_shift_net_x14 <= shift;
  sync_net_x2 <= sync;
  of_x0 <= logical1_y_net_x14;
  pol0_out <= reinterpret1_output_port_net_x4;
  pol1_out <= reinterpret1_output_port_net_x5;
  pol2_out <= reinterpret1_output_port_net_x6;
  pol3_out <= reinterpret1_output_port_net_x7;
  sync_out <= sync_delay1_q_net_x2;

  bi_real_unscr_4x_b9d413eca4: entity work.bi_real_unscr_4x_entity_b9d413eca4
    port map (
      ce_1 => ce_1_sg_x538,
      clk_1 => clk_1_sg_x538,
      even => reinterpret2_output_port_net_x16,
      odd => reinterpret1_output_port_net_x25,
      sync => delay0_q_net_x15,
      pol1_out => reinterpret1_output_port_net_x20,
      pol2_out => reinterpret1_output_port_net_x21,
      pol3_out => reinterpret1_output_port_net_x22,
      pol4_out => reinterpret1_output_port_net_x23,
      sync_out => sync_delay1_q_net_x2
    );

  biplex_core_07162b7c67: entity work.biplex_core_entity_07162b7c67
    port map (
      ce_1 => ce_1_sg_x538,
      clk_1 => clk_1_sg_x538,
      pol1 => reinterpret1_output_port_net_x24,
      pol2 => reinterpret1_output_port_net_x26,
      shift => fft_shift_net_x14,
      sync => sync_net_x2,
      of_x0 => logical1_y_net_x14,
      out1 => reinterpret2_output_port_net_x16,
      out2 => reinterpret1_output_port_net_x25,
      sync_out => delay0_q_net_x15
    );

  even_bussify_62b3b2aba4: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => concat_y_net_x1,
      bus_out => reinterpret1_output_port_net_x24
    );

  odd_bussify_4e0475bdea: entity work.d_bussify_entity_edab46ac75
    port map (
      in1 => concat_y_net_x2,
      bus_out => reinterpret1_output_port_net_x26
    );

  pol0_debus_14d3dd05ce: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x20,
      msb_lsb_out1 => reinterpret1_output_port_net_x4
    );

  pol1_debus_0626428a1c: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x21,
      msb_lsb_out1 => reinterpret1_output_port_net_x5
    );

  pol2_debus_f7e12b655a: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x22,
      msb_lsb_out1 => reinterpret1_output_port_net_x6
    );

  pol3_debus_484c5c53cc: entity work.expand0_entity_49f6172f66
    port map (
      bus_in => reinterpret1_output_port_net_x23,
      msb_lsb_out1 => reinterpret1_output_port_net_x7
    );

  ri_to_c0_ec70da5d21: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => pol2_net_x1,
      re => pol1_net_x1,
      c => concat_y_net_x1
    );

  ri_to_c1_63ae11e57b: entity work.ri_to_c_entity_5ed22bc0d3
    port map (
      im => pol4_net_x1,
      re => pol3_net_x1,
      c => concat_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "fft_astro_devel_core"

entity fft_astro_devel_core is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_shift: in std_logic_vector(31 downto 0); 
    pol1: in std_logic_vector(17 downto 0); 
    pol2: in std_logic_vector(17 downto 0); 
    pol3: in std_logic_vector(17 downto 0); 
    pol4: in std_logic_vector(17 downto 0); 
    sync: in std_logic; 
    fft_oflow: out std_logic; 
    out_pol1: out std_logic_vector(35 downto 0); 
    out_pol2: out std_logic_vector(35 downto 0); 
    out_pol3: out std_logic_vector(35 downto 0); 
    out_pol4: out std_logic_vector(35 downto 0); 
    sync_out: out std_logic
  );
end fft_astro_devel_core;

architecture structural of fft_astro_devel_core is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "fft_astro_devel_core,sysgen_core,{clock_period=10.00000000,clocking=Clock_Enables,compilation=NGC_Netlist,sample_periods=1.00000000000,testbench=0,total_blocks=13236,xilinx_adder_subtracter_block=242,xilinx_arithmetic_relational_operator_block=50,xilinx_assert_block=11,xilinx_bit_slice_extractor_block=1578,xilinx_bus_concatenator_block=461,xilinx_bus_multiplexer_block=134,xilinx_constant_block_block=452,xilinx_counter_block=53,xilinx_delay_block=733,xilinx_dual_port_random_access_memory_block=7,xilinx_gateway_in_block=6,xilinx_gateway_out_block=6,xilinx_input_scaler_block=60,xilinx_inverter_block=148,xilinx_logical_block_block=326,xilinx_multiplier_block=44,xilinx_negate_block_block=27,xilinx_single_port_random_access_memory_block=82,xilinx_single_port_read_only_memory_block=7,xilinx_system_generator_block=1,xilinx_type_converter_block=96,xilinx_type_reinterpreter_block=2434,}";

  signal ce_1_sg_x539: std_logic;
  signal clk_1_sg_x539: std_logic;
  signal fft_oflow_net: std_logic;
  signal fft_shift_net: std_logic_vector(31 downto 0);
  signal out_pol1_net: std_logic_vector(35 downto 0);
  signal out_pol2_net: std_logic_vector(35 downto 0);
  signal out_pol3_net: std_logic_vector(35 downto 0);
  signal out_pol4_net: std_logic_vector(35 downto 0);
  signal pol1_net: std_logic_vector(17 downto 0);
  signal pol2_net: std_logic_vector(17 downto 0);
  signal pol3_net: std_logic_vector(17 downto 0);
  signal pol4_net: std_logic_vector(17 downto 0);
  signal sync_net: std_logic;
  signal sync_out_net: std_logic;

begin
  ce_1_sg_x539 <= ce_1;
  clk_1_sg_x539 <= clk_1;
  fft_shift_net <= fft_shift;
  pol1_net <= pol1;
  pol2_net <= pol2;
  pol3_net <= pol3;
  pol4_net <= pol4;
  sync_net <= sync;
  fft_oflow <= fft_oflow_net;
  out_pol1 <= out_pol1_net;
  out_pol2 <= out_pol2_net;
  out_pol3 <= out_pol3_net;
  out_pol4 <= out_pol4_net;
  sync_out <= sync_out_net;

  fft_biplex_real_4x_f257ec0d37: entity work.fft_biplex_real_4x_entity_f257ec0d37
    port map (
      ce_1 => ce_1_sg_x539,
      clk_1 => clk_1_sg_x539,
      pol0_in => pol1_net,
      pol1_in => pol2_net,
      pol2_in => pol3_net,
      pol3_in => pol4_net,
      shift => fft_shift_net,
      sync => sync_net,
      of_x0 => fft_oflow_net,
      pol0_out => out_pol1_net,
      pol1_out => out_pol2_net,
      pol2_out => out_pol3_net,
      pol3_out => out_pol4_net,
      sync_out => sync_out_net
    );

end structural;
